module epRISC_embeddedROM(iClk, iAddr, oData, iEnable);

    input iClk, iEnable;
    input [11:0] iAddr;
    output wire [31:0] oData;
    
    reg [31:0] rDataOut, rContents[0:4095];
    
    assign oData = (iEnable) ? rDataOut : 32'bz;
    
    always @(posedge iClk) begin
        rDataOut = rContents[iAddr];
    end
    
    initial begin
rContents[0] = 32'h21001100;
rContents[1] = 32'hD0000010;
rContents[2] = 32'h24000007;
rContents[3] = 32'h61400000;
rContents[4] = 32'hD00000CC;
rContents[5] = 32'h41400000;
rContents[6] = 32'h8000011B;
rContents[7] = 32'h65705249;
rContents[8] = 32'h53432042;
rContents[9] = 32'h6F6F746C;
rContents[10] = 32'h6F616465;
rContents[11] = 32'h72207633;
rContents[12] = 32'h202D2073;
rContents[13] = 32'h74617274;
rContents[14] = 32'h696E672E;
rContents[15] = 32'h2E2E0A0D;
rContents[16] = 32'h00000000;
rContents[17] = 32'h61C00000;
rContents[18] = 32'h2C002000;
rContents[19] = 32'h2F010001;
rContents[20] = 32'h6CF00000;
rContents[21] = 32'h04000000;
rContents[22] = 32'h04000000;
rContents[23] = 32'h04000000;
rContents[24] = 32'h04000000;
rContents[25] = 32'h41C00000;
rContents[26] = 32'hF0000000;
rContents[27] = 32'h61E00000;
rContents[28] = 32'h61D00000;
rContents[29] = 32'h61C00000;
rContents[30] = 32'h18111004;
rContents[31] = 32'h2C002000;
rContents[32] = 32'h41D00000;
rContents[33] = 32'h41E00000;
rContents[34] = 32'h2F600008;
rContents[35] = 32'h103FFE00;
rContents[36] = 32'h186FF010;
rContents[37] = 32'h103FFD00;
rContents[38] = 32'h6CF00001;
rContents[39] = 32'h2F010005;
rContents[40] = 32'h6CF00000;
rContents[41] = 32'h4CF00000;
rContents[42] = 32'h18F0F001;
rContents[43] = 32'h820FFFFE;
rContents[44] = 32'h4CF00002;
rContents[45] = 32'h18011006;
rContents[46] = 32'h41C00000;
rContents[47] = 32'h41D00000;
rContents[48] = 32'h41E00000;
rContents[49] = 32'hF0000000;
rContents[50] = 32'h61E00000;
rContents[51] = 32'h61C00000;
rContents[52] = 32'h18111003;
rContents[53] = 32'h2C002000;
rContents[54] = 32'h41E00000;
rContents[55] = 32'h2F600000;
rContents[56] = 32'h103FFE00;
rContents[57] = 32'h186FF010;
rContents[58] = 32'h6CF00001;
rContents[59] = 32'h2F010005;
rContents[60] = 32'h6CF00000;
rContents[61] = 32'h4CF00000;
rContents[62] = 32'h18F0F001;
rContents[63] = 32'h820FFFFE;
rContents[64] = 32'h2F600000;
rContents[65] = 32'h103FFE00;
rContents[66] = 32'h186FF010;
rContents[67] = 32'h6CF00001;
rContents[68] = 32'h2F010005;
rContents[69] = 32'h6CF00000;
rContents[70] = 32'h4CF00000;
rContents[71] = 32'h18F0F001;
rContents[72] = 32'h820FFFFE;
rContents[73] = 32'h4CF00002;
rContents[74] = 32'h18011004;
rContents[75] = 32'h41C00000;
rContents[76] = 32'h41E00000;
rContents[77] = 32'hF0000000;
rContents[78] = 32'h61D00000;
rContents[79] = 32'h61C00000;
rContents[80] = 32'h18111003;
rContents[81] = 32'h2C002000;
rContents[82] = 32'h41D00000;
rContents[83] = 32'h2F800100;
rContents[84] = 32'h6CF00001;
rContents[85] = 32'h2F010005;
rContents[86] = 32'h6CF00000;
rContents[87] = 32'h4CF00000;
rContents[88] = 32'h18F0F001;
rContents[89] = 32'h820FFFFE;
rContents[90] = 32'h2F800100;
rContents[91] = 32'h6CF00001;
rContents[92] = 32'h2F010005;
rContents[93] = 32'h6CF00000;
rContents[94] = 32'h4CF00000;
rContents[95] = 32'h18F0F001;
rContents[96] = 32'h820FFFFE;
rContents[97] = 32'h4CF00002;
rContents[98] = 32'h18F0F080;
rContents[99] = 32'h820FFFF7;
rContents[100] = 32'h2F808101;
rContents[101] = 32'h103FFD00;
rContents[102] = 32'h6CF00001;
rContents[103] = 32'h2F010005;
rContents[104] = 32'h6CF00000;
rContents[105] = 32'h4CF00000;
rContents[106] = 32'h18F0F001;
rContents[107] = 32'h820FFFFE;
rContents[108] = 32'h2F808100;
rContents[109] = 32'h3F000080;
rContents[110] = 32'h6CF00001;
rContents[111] = 32'h2F010005;
rContents[112] = 32'h6CF00000;
rContents[113] = 32'h4CF00000;
rContents[114] = 32'h18F0F001;
rContents[115] = 32'h820FFFFE;
rContents[116] = 32'h18011004;
rContents[117] = 32'h41C00000;
rContents[118] = 32'h41D00000;
rContents[119] = 32'hF0000000;
rContents[120] = 32'h61C00000;
rContents[121] = 32'h2C002000;
rContents[122] = 32'h2F808100;
rContents[123] = 32'h3F000020;
rContents[124] = 32'h6CF00001;
rContents[125] = 32'h2F010005;
rContents[126] = 32'h6CF00000;
rContents[127] = 32'h4CF00000;
rContents[128] = 32'h18F0F001;
rContents[129] = 32'h820FFFFE;
rContents[130] = 32'h2F800100;
rContents[131] = 32'h6CF00001;
rContents[132] = 32'h2F010005;
rContents[133] = 32'h6CF00000;
rContents[134] = 32'h4CF00000;
rContents[135] = 32'h18F0F001;
rContents[136] = 32'h820FFFFE;
rContents[137] = 32'h2F800100;
rContents[138] = 32'h6CF00001;
rContents[139] = 32'h2F010005;
rContents[140] = 32'h6CF00000;
rContents[141] = 32'h4CF00000;
rContents[142] = 32'h18F0F001;
rContents[143] = 32'h820FFFFE;
rContents[144] = 32'h4CF00002;
rContents[145] = 32'h18F0F020;
rContents[146] = 32'h820FFFF7;
rContents[147] = 32'h2F800102;
rContents[148] = 32'h6CF00001;
rContents[149] = 32'h2F010005;
rContents[150] = 32'h6CF00000;
rContents[151] = 32'h4CF00000;
rContents[152] = 32'h18F0F001;
rContents[153] = 32'h820FFFFE;
rContents[154] = 32'h2F800102;
rContents[155] = 32'h6CF00001;
rContents[156] = 32'h2F010005;
rContents[157] = 32'h6CF00000;
rContents[158] = 32'h4CF00000;
rContents[159] = 32'h18F0F001;
rContents[160] = 32'h820FFFFE;
rContents[161] = 32'h4CF00002;
rContents[162] = 32'h41C00000;
rContents[163] = 32'hF0000000;
rContents[164] = 32'h61C00000;
rContents[165] = 32'h61D00000;
rContents[166] = 32'h61E00000;
rContents[167] = 32'h18111004;
rContents[168] = 32'h41C00000;
rContents[169] = 32'h2E000008;
rContents[170] = 32'h18011005;
rContents[171] = 32'h182DCCF0;
rContents[172] = 32'h186CC004;
rContents[173] = 32'h188DD01C;
rContents[174] = 32'h180DD030;
rContents[175] = 32'h18E0D03A;
rContents[176] = 32'h83000002;
rContents[177] = 32'h180DD007;
rContents[178] = 32'h61D00000;
rContents[179] = 32'hD00FFF9B;
rContents[180] = 32'h41D00000;
rContents[181] = 32'h181EE001;
rContents[182] = 32'h18E0E000;
rContents[183] = 32'h8D0FFFF4;
rContents[184] = 32'h41E00000;
rContents[185] = 32'h41D00000;
rContents[186] = 32'h41C00000;
rContents[187] = 32'hF0000000;
rContents[188] = 32'h61C00000;
rContents[189] = 32'h61D00000;
rContents[190] = 32'h61E00000;
rContents[191] = 32'h18111004;
rContents[192] = 32'h41D00000;
rContents[193] = 32'h41C00000;
rContents[194] = 32'h18011006;
rContents[195] = 32'h08ED0000;
rContents[196] = 32'h187DD002;
rContents[197] = 32'h100CCD00;
rContents[198] = 32'h4CF00000;
rContents[199] = 32'h2D000003;
rContents[200] = 32'h182EE003;
rContents[201] = 32'h101EDE00;
rContents[202] = 32'h186EE003;
rContents[203] = 32'h10DFFEFF;
rContents[204] = 32'h41E00000;
rContents[205] = 32'h41D00000;
rContents[206] = 32'h41C00000;
rContents[207] = 32'hF0000000;
rContents[208] = 32'h61C00000;
rContents[209] = 32'h61D00000;
rContents[210] = 32'h18111003;
rContents[211] = 32'h2D000000;
rContents[212] = 32'h41C00000;
rContents[213] = 32'h18011004;
rContents[214] = 32'h61C00000;
rContents[215] = 32'h61D00000;
rContents[216] = 32'hD00FFFE4;
rContents[217] = 32'h41D00000;
rContents[218] = 32'h18E0F000;
rContents[219] = 32'h81000006;
rContents[220] = 32'h61F00000;
rContents[221] = 32'hD00FFF71;
rContents[222] = 32'h41F00000;
rContents[223] = 32'h180DD001;
rContents[224] = 32'h800FFFF7;
rContents[225] = 32'h41C00000;
rContents[226] = 32'h41D00000;
rContents[227] = 32'h41C00000;
rContents[228] = 32'hF0000000;
rContents[229] = 32'h0A0A416E;
rContents[230] = 32'h20657272;
rContents[231] = 32'h6F722068;
rContents[232] = 32'h6173206F;
rContents[233] = 32'h63637572;
rContents[234] = 32'h65642E0A;
rContents[235] = 32'h00000000;
rContents[236] = 32'h0A0A4120;
rContents[237] = 32'h66617461;
rContents[238] = 32'h6C206572;
rContents[239] = 32'h726F7220;
rContents[240] = 32'h68617320;
rContents[241] = 32'h6F636375;
rContents[242] = 32'h7265642E;
rContents[243] = 32'h0A000000;
rContents[244] = 32'h43616C6C;
rContents[245] = 32'h65642061;
rContents[246] = 32'h74200000;
rContents[247] = 32'h53746163;
rContents[248] = 32'h6B747261;
rContents[249] = 32'h63652028;
rContents[250] = 32'h746F7020;
rContents[251] = 32'h3136293A;
rContents[252] = 32'h0A000000;
rContents[253] = 32'h52656769;
rContents[254] = 32'h73746572;
rContents[255] = 32'h733A0A00;
rContents[256] = 32'h52657375;
rContents[257] = 32'h6D696E67;
rContents[258] = 32'h2E0A0A00;
rContents[259] = 32'h48616C74;
rContents[260] = 32'h696E672E;
rContents[261] = 32'h0A0A0000;
rContents[262] = 32'h80000001;
rContents[263] = 32'h2F0000EC;
rContents[264] = 32'h61F00000;
rContents[265] = 32'hD00FFFC7;
rContents[266] = 32'h41F00000;
rContents[267] = 32'h2F0000F4;
rContents[268] = 32'h61F00000;
rContents[269] = 32'hD00FFFC3;
rContents[270] = 32'h41F00000;
rContents[271] = 32'hD00FFF95;
rContents[272] = 32'h04200000;
rContents[273] = 32'hF0000000;
rContents[274] = 32'hF0000000;
rContents[275] = 32'h4C656D6F;
rContents[276] = 32'h6E207630;
rContents[277] = 32'h2E32202D;
rContents[278] = 32'h20666F72;
rContents[279] = 32'h20657052;
rContents[280] = 32'h49534320;
rContents[281] = 32'h76352073;
rContents[282] = 32'h79737465;
rContents[283] = 32'h6D730000;
rContents[284] = 32'h800FFF32;
rContents[285] = 32'h800FFF5B;
rContents[286] = 32'h800FFF86;
rContents[287] = 32'h800FFFB1;
rContents[288] = 32'h800FFFE7;
rContents[289] = 32'h210017FF;
rContents[290] = 32'h28000113;
rContents[291] = 32'h61800000;
rContents[292] = 32'hD00FFFFB;
rContents[293] = 32'h41800000;
rContents[294] = 32'h26001000;
rContents[295] = 32'h29000000;
rContents[296] = 32'h2800000A;
rContents[297] = 32'h61800000;
rContents[298] = 32'hD00FFFF2;
rContents[299] = 32'h41800000;
rContents[300] = 32'h2800000D;
rContents[301] = 32'h61800000;
rContents[302] = 32'hD00FFFEE;
rContents[303] = 32'h41800000;
rContents[304] = 32'h2800003E;
rContents[305] = 32'h61800000;
rContents[306] = 32'hD00FFFEA;
rContents[307] = 32'h41800000;
rContents[308] = 32'hD00FFFE9;
rContents[309] = 32'h18E0F008;
rContents[310] = 32'h82000008;
rContents[311] = 32'h18166001;
rContents[312] = 32'h18199001;
rContents[313] = 32'h46F00000;
rContents[314] = 32'h61F00000;
rContents[315] = 32'hD00FFFE1;
rContents[316] = 32'h41F00000;
rContents[317] = 32'h800FFFF7;
rContents[318] = 32'h18E0F00D;
rContents[319] = 32'h82000003;
rContents[320] = 32'h66F00000;
rContents[321] = 32'h8000000A;
rContents[322] = 32'h18F09180;
rContents[323] = 32'h820FFFF1;
rContents[324] = 32'h61F00000;
rContents[325] = 32'hD00FFFD7;
rContents[326] = 32'h41F00000;
rContents[327] = 32'h66F00000;
rContents[328] = 32'h18066001;
rContents[329] = 32'h18099001;
rContents[330] = 32'h800FFFEA;
rContents[331] = 32'h26001000;
rContents[332] = 32'h2800000A;
rContents[333] = 32'h61800000;
rContents[334] = 32'hD00FFFCE;
rContents[335] = 32'h41800000;
rContents[336] = 32'h2800000D;
rContents[337] = 32'h61800000;
rContents[338] = 32'hD00FFFCA;
rContents[339] = 32'h41800000;
rContents[340] = 32'h46900000;
rContents[341] = 32'h18E0900D;
rContents[342] = 32'h82000005;
rContents[343] = 32'h18E0703A;
rContents[344] = 32'h82000002;
rContents[345] = 32'h41800000;
rContents[346] = 32'h800FFFCC;
rContents[347] = 32'h18E09052;
rContents[348] = 32'h82000003;
rContents[349] = 32'hD0400000;
rContents[350] = 32'h800FFFF6;
rContents[351] = 32'h18E0903A;
rContents[352] = 32'h82000005;
rContents[353] = 32'h2700003A;
rContents[354] = 32'h61400000;
rContents[355] = 32'h18066001;
rContents[356] = 32'h800FFFF0;
rContents[357] = 32'h18E0902E;
rContents[358] = 32'h82000007;
rContents[359] = 32'h18E0703A;
rContents[360] = 32'h82000002;
rContents[361] = 32'h41800000;
rContents[362] = 32'h2700002E;
rContents[363] = 32'h18066001;
rContents[364] = 32'h800FFFE8;
rContents[365] = 32'h18E09020;
rContents[366] = 32'h82000003;
rContents[367] = 32'h18066001;
rContents[368] = 32'h800FFFE4;
rContents[369] = 32'h25000000;
rContents[370] = 32'h46900000;
rContents[371] = 32'h18199030;
rContents[372] = 32'h18E0900A;
rContents[373] = 32'h84000005;
rContents[374] = 32'h18199007;
rContents[375] = 32'h18E09010;
rContents[376] = 32'h84000002;
rContents[377] = 32'h80000005;
rContents[378] = 32'h18655004;
rContents[379] = 32'h10355900;
rContents[380] = 32'h18066001;
rContents[381] = 32'h800FFFF5;
rContents[382] = 32'h46900000;
rContents[383] = 32'h18E0703A;
rContents[384] = 32'h82000004;
rContents[385] = 32'h64500000;
rContents[386] = 32'h18044001;
rContents[387] = 32'h800FFFD1;
rContents[388] = 32'h61400000;
rContents[389] = 32'h08450000;
rContents[390] = 32'h18E0703A;
rContents[391] = 32'h82000003;
rContents[392] = 32'h41800000;
rContents[393] = 32'h800FFFCB;
rContents[394] = 32'h18E0703A;
rContents[395] = 32'h8200001A;
rContents[396] = 32'h41800000;
rContents[397] = 32'h61400000;
rContents[398] = 32'hD00FFF16;
rContents[399] = 32'h41400000;
rContents[400] = 32'h2800003E;
rContents[401] = 32'h61800000;
rContents[402] = 32'hD00FFF8A;
rContents[403] = 32'h41800000;
rContents[404] = 32'h28000020;
rContents[405] = 32'h61800000;
rContents[406] = 32'hD00FFF86;
rContents[407] = 32'h41800000;
rContents[408] = 32'h44800000;
rContents[409] = 32'h61800000;
rContents[410] = 32'hD00FFF84;
rContents[411] = 32'h41400000;
rContents[412] = 32'h2800000A;
rContents[413] = 32'h61800000;
rContents[414] = 32'hD00FFF7E;
rContents[415] = 32'h41800000;
rContents[416] = 32'h2800000D;
rContents[417] = 32'h61800000;
rContents[418] = 32'hD00FFF7A;
rContents[419] = 32'h41800000;
rContents[420] = 32'h800FFFB0;
rContents[421] = 32'h18E0703A;
rContents[422] = 32'hD20FFF7A;
rContents[423] = 32'h08840000;
rContents[424] = 32'h41400000;
rContents[425] = 32'h101A8400;
rContents[426] = 32'h80000009;
rContents[427] = 32'h2800000A;
rContents[428] = 32'h61800000;
rContents[429] = 32'hD00FFF6F;
rContents[430] = 32'h41800000;
rContents[431] = 32'h2800000D;
rContents[432] = 32'h61800000;
rContents[433] = 32'hD00FFF6B;
rContents[434] = 32'h41800000;
rContents[435] = 32'h61400000;
rContents[436] = 32'hD00FFEF0;
rContents[437] = 32'h41400000;
rContents[438] = 32'h2800003E;
rContents[439] = 32'h61800000;
rContents[440] = 32'hD00FFF64;
rContents[441] = 32'h41800000;
rContents[442] = 32'h18E0A007;
rContents[443] = 32'h89000003;
rContents[444] = 32'h08BA0000;
rContents[445] = 32'h80000002;
rContents[446] = 32'h2B000008;
rContents[447] = 32'h101AAB00;
rContents[448] = 32'h28000020;
rContents[449] = 32'h61800000;
rContents[450] = 32'hD00FFF5A;
rContents[451] = 32'h41800000;
rContents[452] = 32'h44800000;
rContents[453] = 32'h61800000;
rContents[454] = 32'hD00FFF58;
rContents[455] = 32'h41400000;
rContents[456] = 32'h18044001;
rContents[457] = 32'h181BB001;
rContents[458] = 32'h18E0B000;
rContents[459] = 32'h810FFFF5;
rContents[460] = 32'h18E0A000;
rContents[461] = 32'h820FFFDE;
rContents[462] = 32'h800FFF86;
    end

endmodule

/*  Program 1 - square wave generator over GPIO
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808000;
        rContents[8] = 32'h3500FFFF;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25000000;
        rContents[17] = 32'h08650000;
        rContents[18] = 32'h36808002;
        rContents[19] = 32'h64600001;
        rContents[20] = 32'h27010005;
        rContents[21] = 32'h64700000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h04000000;
        rContents[26] = 32'h18B5580F;
        rContents[27] = 32'h18055001;
        rContents[28] = 32'h800FFFF5;
        rContents[29] = 32'h0;
        rContents[30] = 32'h0;
        rContents[31] = 32'h0;
        rContents[32] = 32'h0;
        rContents[33] = 32'h0;
        rContents[34] = 32'h0;
        rContents[35] = 32'h0; */
        
/*  Program 2 - print some 'H's over the serial link
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808101;
        rContents[8] = 32'h35000048;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25808100;
        rContents[17] = 32'h35000080;
        rContents[18] = 32'h64500001;
        rContents[19] = 32'h27010005;
        rContents[20] = 32'h64700000;
        rContents[21] = 32'h04000000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h800FFFED; */
