/* verilator lint_off WIDTH */

module epRISC_VideoTerm(iClk, iRst, iAddr, iData, oData, iWrite, iEnable, iMemClk, iVideoClk, oColor, oHS, oVS);

    input iClk, iRst, iWrite, iEnable, iMemClk, iVideoClk;
    input [1:0] iAddr;
    input [15:0] iData;
    output wire [7:0] oColor;
    output reg oHS, oVS;
    output wire [15:0] oData;
    
    reg [3:0] rRowSel;
    reg [7:0] rDataOutput, rColorOutput;
    reg [9:0] rPulseX, rPulseY;
    reg [11:0] rTempX, rTempY, rFramePtr;
    reg [15:0] rConfig, rRow, rColumn;
    
    wire mDrawingValidLine, mDrawingValidFrame, mDrawingValidData;
    wire [7:0] wCurrColor, wCurrChar, wFontRow;
    wire [9:0] wPixelX, wPixelY;
    wire [15:0] wCharRAMData, wCharRAMFrame;
        
    assign oData = (!iEnable) ? 16'bz : ((iAddr==0)?rConfig:((iAddr==1)?rColumn:((iAddr==2)?rRow:((iAddr==3)?wCharRAMData:16'b1))));
    
    assign oColor = (rDataOutput[7-wPixelX[2:0]] && mDrawingValidData) ? rColorOutput : 8'h0; //either color or black
    //(mDrawingValidData && ((wPixelX[0] && wPixelY[0]) || (!wPixelX[0] && !wPixelY[0]))) ? 8'hFF : 8'h0; //this is a fine-checkerboard test pattern

    assign mDrawingValidLine = (rPulseY >= 35 && rPulseY < 515) ? 1 : 0;
    assign mDrawingValidFrame = (rPulseX >= 160 && rPulseX < 800) ? 1 : 0;
    assign mDrawingValidData = (mDrawingValidLine && mDrawingValidFrame) ? 1 : 0;
    
    assign wPixelX = rPulseX - 10'd160;
    assign wPixelY = rPulseY - 10'd35;
       
    assign wCurrColor = wCharRAMFrame[15:8];
    assign wCurrChar = wCharRAMFrame[7:0];
    
    wire [16:0] debug;
    assign debug = (rRow<<4)+(rRow<<6)+rColumn;
    
    `ifdef EMULATED
    SoftVideoRAM vram((rRow<<4)+(rRow<<6)+rColumn, rFramePtr[11:0], iClk, iMemClk, iData, 16'h0, (iWrite&&iEnable&&iAddr==3)?1:0, 0, wCharRAMData, wCharRAMFrame);
    `else
    ChipVideoRAM vram((rRow<<4)+(rRow<<6)+rColumn, rFramePtr[11:0], iClk, iMemClk, iData, 16'h0, (iWrite&&iEnable&&iAddr==3)?1:0, 0, wCharRAMData, wCharRAMFrame);
    `endif
    
    VideoROM vrom({rRowSel, wCurrChar}, iMemClk, wFontRow);
    
    always @(posedge iClk) begin
        if(iRst) begin
            rConfig <= 16'h0;
        end else begin
            if(iWrite && iEnable && (iAddr == 0))
                rConfig <= iData;
        end
    end

    always @(posedge iClk) begin
        if(iRst) begin
            rRow <= 16'h0;
        end else begin
            if(iWrite && iEnable && (iAddr == 2))
                rRow <= iData;
        end
    end
    
    always @(posedge iClk) begin
        if(iRst) begin
            rColumn <= 16'h0;
        end else begin
            if(iWrite && iEnable && (iAddr == 1))
                rColumn <= iData;
        end
    end
        
    always @(posedge iVideoClk) begin
        if(iRst) begin
            rPulseX <= 0;
            rPulseY <= 0;
            rRowSel <= 0;
        end else begin
            rPulseX <= rPulseX + 1;
            
            case(rPulseX)
                0: oHS <= 1;
                16: oHS <= 0;
                112: oHS <= 1;
                800: begin rPulseY <= rPulseY + 1; rRowSel <= rRowSel + 1; rPulseX <= 0; end
            endcase
            
            case(rPulseY)
                0: oVS <= 1;
                10: oVS <= 0;
                12: oVS <= 1;
                525: begin rPulseY <= 0; rRowSel <= 0; end
            endcase
            
            if(rRowSel == 12)
                rRowSel <= 0;
        end
    end

    always @(posedge iVideoClk) begin
        if(iRst) begin
            rDataOutput <= 0;
            rFramePtr <= 0;
        end else begin
            //rFramePtr <= 0;
            
            case(wPixelX[2:0])
                3'h6: begin
                    if(rPulseX < 154) begin
                        rTempX <= 0;
                    end else if(rPulseX >= 154 && rPulseX < 160) begin
                        rTempX <= 1;
                    end else begin
                        rTempX <= 2 + (wPixelX / 8);
                    end
                    
                    rTempY <= wPixelY / 12;
                    rFramePtr <= (rTempY * 80) + rTempX;
                end
                
                3'h7: begin
                    rDataOutput <= wFontRow;
                    rColorOutput <= wCurrColor;
                end
            endcase
        end
    end
    
endmodule

module SoftVideoRAM(iAddrA, iAddrB, iClkA, iClkB, iDInA, iDInB, iWriteA, iWriteB, oDOutA, oDOutB);
    input iClkA, iClkB, iWriteA, iWriteB;
    input [11:0] iAddrA, iAddrB;
    input [15:0] iDInA, iDInB;
    output reg [15:0] oDOutA, oDOutB;
    
    reg [12:0] rClr;
    reg [15:0] rContents[0:4095];

    wire debug;
    assign debug = (iAddrB > 80) ? 1 : 0;
    
    initial begin
        for(rClr=0;rClr<4096;rClr=rClr+1)
            rContents[rClr] = 0;
    end
    
    always @(posedge iClkA) begin
        if(iWriteA) begin
            rContents[iAddrA] <= iDInA;
        end
    end
    
    always @(posedge iClkB) begin
        if(iWriteB) begin
            rContents[iAddrB] <= iDInB;
        end
    end
    
    always @(posedge iClkA) begin
        if(!iWriteA) begin
            oDOutA <= rContents[iAddrA];
        end
    end
    
    always @(posedge iClkB) begin
        if(!iWriteB) begin
            oDOutB <= rContents[iAddrB];
        end
    end
endmodule

module VideoROM(iAddr, iClk, oData);

    input iClk;
    input [11:0] iAddr;
    output wire [15:0] oData;
    
    reg [15:0] rDataOut, rContents[0:3071];
    
    assign oData = rDataOut;
    
    always @(posedge iClk) begin
        rDataOut = rContents[iAddr];
    end
    
    initial begin
        rContents[0] = 8'b01010101;
        rContents[1] = 8'b10101010;
        rContents[2] = 8'b01010101;
        rContents[3] = 8'b11111111;
        rContents[4] = 8'b11111111;
        rContents[5] = 8'b00000000;
        rContents[6] = 8'b11111110;
        rContents[7] = 8'b11111110;
        rContents[8] = 8'b00111000;
        rContents[9] = 8'b01111100;
        rContents[10] = 8'b01111100;
        rContents[11] = 8'b01101100;
        rContents[12] = 8'b00010000;
        rContents[13] = 8'b00111000;
        rContents[14] = 8'b00010000;
        rContents[15] = 8'b11111110;
        rContents[16] = 8'b11111110;
        rContents[17] = 8'b11111110;
        rContents[18] = 8'b00111000;
        rContents[19] = 8'b00111110;
        rContents[20] = 8'b00010000;
        rContents[21] = 8'b00010000;
        rContents[22] = 8'b00000000;
        rContents[23] = 8'b00000000;
        rContents[24] = 8'b11000000;
        rContents[25] = 8'b00000110;
        rContents[26] = 8'b00010000;
        rContents[27] = 8'b11111110;
        rContents[28] = 8'b00010000;
        rContents[29] = 8'b00000000;
        rContents[30] = 8'b00010000;
        rContents[31] = 8'b01111100;
        rContents[32] = 8'b00000000;
        rContents[33] = 8'b00010000;
        rContents[34] = 8'b00101000;
        rContents[35] = 8'b01000100;
        rContents[36] = 8'b00010000;
        rContents[37] = 8'b11100010;
        rContents[38] = 8'b11111110;
        rContents[39] = 8'b00010000;
        rContents[40] = 8'b00001000;
        rContents[41] = 8'b00100000;
        rContents[42] = 8'b00010000;
        rContents[43] = 8'b00000000;
        rContents[44] = 8'b00000000;
        rContents[45] = 8'b00000000;
        rContents[46] = 8'b00000000;
        rContents[47] = 8'b00000010;
        rContents[48] = 8'b01111100;
        rContents[49] = 8'b00010000;
        rContents[50] = 8'b01111100;
        rContents[51] = 8'b01111100;
        rContents[52] = 8'b10000010;
        rContents[53] = 8'b11111110;
        rContents[54] = 8'b01111110;
        rContents[55] = 8'b11111110;
        rContents[56] = 8'b01111100;
        rContents[57] = 8'b01111100;
        rContents[58] = 8'b00000000;
        rContents[59] = 8'b00000000;
        rContents[60] = 8'b00000010;
        rContents[61] = 8'b00000000;
        rContents[62] = 8'b10000000;
        rContents[63] = 8'b01111100;
        rContents[64] = 8'b11111100;
        rContents[65] = 8'b00000110;
        rContents[66] = 8'b11111110;
        rContents[67] = 8'b11111110;
        rContents[68] = 8'b11111100;
        rContents[69] = 8'b11111110;
        rContents[70] = 8'b11111110;
        rContents[71] = 8'b11111110;
        rContents[72] = 8'b10000010;
        rContents[73] = 8'b11111110;
        rContents[74] = 8'b00000010;
        rContents[75] = 8'b10000010;
        rContents[76] = 8'b10000000;
        rContents[77] = 8'b11111110;
        rContents[78] = 8'b10000010;
        rContents[79] = 8'b11111110;
        rContents[80] = 8'b11111110;
        rContents[81] = 8'b11111110;
        rContents[82] = 8'b11111110;
        rContents[83] = 8'b11111110;
        rContents[84] = 8'b11111110;
        rContents[85] = 8'b10000010;
        rContents[86] = 8'b10000010;
        rContents[87] = 8'b10000010;
        rContents[88] = 8'b10000010;
        rContents[89] = 8'b10000010;
        rContents[90] = 8'b11111110;
        rContents[91] = 8'b00111000;
        rContents[92] = 8'b10000000;
        rContents[93] = 8'b00111000;
        rContents[94] = 8'b00010000;
        rContents[95] = 8'b00000000;
        rContents[96] = 8'b00100000;
        rContents[97] = 8'b00000000;
        rContents[98] = 8'b10000000;
        rContents[99] = 8'b00000000;
        rContents[100] = 8'b00000010;
        rContents[101] = 8'b00000000;
        rContents[102] = 8'b11111110;
        rContents[103] = 8'b00000000;
        rContents[104] = 8'b10000000;
        rContents[105] = 8'b00000000;
        rContents[106] = 8'b00000000;
        rContents[107] = 8'b10000000;
        rContents[108] = 8'b00010000;
        rContents[109] = 8'b00000000;
        rContents[110] = 8'b00000000;
        rContents[111] = 8'b00000000;
        rContents[112] = 8'b00000000;
        rContents[113] = 8'b00000000;
        rContents[114] = 8'b00000000;
        rContents[115] = 8'b00000000;
        rContents[116] = 8'b10000000;
        rContents[117] = 8'b00000000;
        rContents[118] = 8'b00000000;
        rContents[119] = 8'b00000000;
        rContents[120] = 8'b00000000;
        rContents[121] = 8'b00000000;
        rContents[122] = 8'b00000000;
        rContents[123] = 8'b00011000;
        rContents[124] = 8'b00010000;
        rContents[125] = 8'b00110000;
        rContents[126] = 8'b00000000;
        rContents[127] = 8'b00010000;
        rContents[128] = 8'b00010000;
        rContents[129] = 8'b11111111;
        rContents[130] = 8'b11111111;
        rContents[131] = 8'b11110000;
        rContents[132] = 8'b00001111;
        rContents[133] = 8'b11110000;
        rContents[134] = 8'b00001111;
        rContents[135] = 8'b00000000;
        rContents[136] = 8'b00000000;
        rContents[137] = 8'b11110000;
        rContents[138] = 8'b00001111;
        rContents[139] = 8'b11111111;
        rContents[140] = 8'b00000000;
        rContents[141] = 8'b00011000;
        rContents[142] = 8'b00000000;
        rContents[143] = 8'b00011000;
        rContents[144] = 8'b00011000;
        rContents[145] = 8'b00000000;
        rContents[146] = 8'b00000000;
        rContents[147] = 8'b00011000;
        rContents[148] = 8'b00000000;
        rContents[149] = 8'b00011000;
        rContents[150] = 8'b00011000;
        rContents[151] = 8'b00011000;
        rContents[152] = 8'b00100100;
        rContents[153] = 8'b00000000;
        rContents[154] = 8'b00100100;
        rContents[155] = 8'b00100100;
        rContents[156] = 8'b00000000;
        rContents[157] = 8'b00000000;
        rContents[158] = 8'b00100100;
        rContents[159] = 8'b00000000;
        rContents[160] = 8'b00100100;
        rContents[161] = 8'b00100100;
        rContents[162] = 8'b00111000;
        rContents[163] = 8'b00000000;
        rContents[164] = 8'b00000000;
        rContents[165] = 8'b11111100;
        rContents[166] = 8'b11111110;
        rContents[167] = 8'b00000110;
        rContents[168] = 8'b00000000;
        rContents[169] = 8'b00000000;
        rContents[170] = 8'b00000000;
        rContents[171] = 8'b00000000;
        rContents[172] = 8'b00000000;
        rContents[173] = 8'b00000000;
        rContents[174] = 8'b00000000;
        rContents[175] = 8'b00000000;
        rContents[176] = 8'b00000000;
        rContents[177] = 8'b00000000;
        rContents[178] = 8'b00000000;
        rContents[179] = 8'b00000000;
        rContents[180] = 8'b00000000;
        rContents[181] = 8'b00000000;
        rContents[182] = 8'b00000000;
        rContents[183] = 8'b00000000;
        rContents[184] = 8'b00000000;
        rContents[185] = 8'b00000000;
        rContents[186] = 8'b00000000;
        rContents[187] = 8'b00000000;
        rContents[188] = 8'b00000000;
        rContents[189] = 8'b00000000;
        rContents[190] = 8'b00000000;
        rContents[191] = 8'b00000000;
        rContents[192] = 8'b00000000;
        rContents[193] = 8'b00000000;
        rContents[194] = 8'b00000000;
        rContents[195] = 8'b00000000;
        rContents[196] = 8'b00000000;
        rContents[197] = 8'b00000000;
        rContents[198] = 8'b00000000;
        rContents[199] = 8'b00000000;
        rContents[200] = 8'b00000000;
        rContents[201] = 8'b00000000;
        rContents[202] = 8'b00000000;
        rContents[203] = 8'b00000000;
        rContents[204] = 8'b00000000;
        rContents[205] = 8'b00000000;
        rContents[206] = 8'b00000000;
        rContents[207] = 8'b00000000;
        rContents[208] = 8'b00000000;
        rContents[209] = 8'b00000000;
        rContents[210] = 8'b00000000;
        rContents[211] = 8'b00000000;
        rContents[212] = 8'b00000000;
        rContents[213] = 8'b00000000;
        rContents[214] = 8'b00000000;
        rContents[215] = 8'b00000000;
        rContents[216] = 8'b00000000;
        rContents[217] = 8'b00000000;
        rContents[218] = 8'b00000000;
        rContents[219] = 8'b00000000;
        rContents[220] = 8'b00000000;
        rContents[221] = 8'b00000000;
        rContents[222] = 8'b00000000;
        rContents[223] = 8'b00000000;
        rContents[224] = 8'b00000000;
        rContents[225] = 8'b00000000;
        rContents[226] = 8'b00000000;
        rContents[227] = 8'b00000000;
        rContents[228] = 8'b00000000;
        rContents[229] = 8'b00000000;
        rContents[230] = 8'b00000000;
        rContents[231] = 8'b00000000;
        rContents[232] = 8'b00000000;
        rContents[233] = 8'b00000000;
        rContents[234] = 8'b00000000;
        rContents[235] = 8'b00000000;
        rContents[236] = 8'b00000000;
        rContents[237] = 8'b00000000;
        rContents[238] = 8'b00000000;
        rContents[239] = 8'b00000000;
        rContents[240] = 8'b00000000;
        rContents[241] = 8'b00000000;
        rContents[242] = 8'b00000000;
        rContents[243] = 8'b00000000;
        rContents[244] = 8'b00000000;
        rContents[245] = 8'b00000000;
        rContents[246] = 8'b00000000;
        rContents[247] = 8'b00000000;
        rContents[248] = 8'b00000000;
        rContents[249] = 8'b00000000;
        rContents[250] = 8'b00000000;
        rContents[251] = 8'b00000000;
        rContents[252] = 8'b00000000;
        rContents[253] = 8'b00000000;
        rContents[254] = 8'b00000000;
        rContents[255] = 8'b00000000;
        rContents[256] = 8'b01010101;
        rContents[257] = 8'b10101010;
        rContents[258] = 8'b11111111;
        rContents[259] = 8'b10101010;
        rContents[260] = 8'b11111111;
        rContents[261] = 8'b00000000;
        rContents[262] = 8'b11111110;
        rContents[263] = 8'b10000010;
        rContents[264] = 8'b00010000;
        rContents[265] = 8'b10000010;
        rContents[266] = 8'b11111110;
        rContents[267] = 8'b11111110;
        rContents[268] = 8'b00111000;
        rContents[269] = 8'b01111100;
        rContents[270] = 8'b00010000;
        rContents[271] = 8'b10000010;
        rContents[272] = 8'b10000010;
        rContents[273] = 8'b11111110;
        rContents[274] = 8'b00100000;
        rContents[275] = 8'b00100010;
        rContents[276] = 8'b00111000;
        rContents[277] = 8'b00010000;
        rContents[278] = 8'b00000000;
        rContents[279] = 8'b00000000;
        rContents[280] = 8'b11110000;
        rContents[281] = 8'b00011110;
        rContents[282] = 8'b00111000;
        rContents[283] = 8'b10001010;
        rContents[284] = 8'b00111000;
        rContents[285] = 8'b00000000;
        rContents[286] = 8'b00111000;
        rContents[287] = 8'b01000000;
        rContents[288] = 8'b00000000;
        rContents[289] = 8'b00010000;
        rContents[290] = 8'b00101000;
        rContents[291] = 8'b01000100;
        rContents[292] = 8'b11111110;
        rContents[293] = 8'b10100010;
        rContents[294] = 8'b10000010;
        rContents[295] = 8'b00010000;
        rContents[296] = 8'b00010000;
        rContents[297] = 8'b00010000;
        rContents[298] = 8'b00101000;
        rContents[299] = 8'b00000000;
        rContents[300] = 8'b00000000;
        rContents[301] = 8'b00000000;
        rContents[302] = 8'b00000000;
        rContents[303] = 8'b00000010;
        rContents[304] = 8'b10000010;
        rContents[305] = 8'b00110000;
        rContents[306] = 8'b10000010;
        rContents[307] = 8'b10000010;
        rContents[308] = 8'b10000010;
        rContents[309] = 8'b10000000;
        rContents[310] = 8'b10000000;
        rContents[311] = 8'b00000010;
        rContents[312] = 8'b10000010;
        rContents[313] = 8'b10000010;
        rContents[314] = 8'b00010000;
        rContents[315] = 8'b00010000;
        rContents[316] = 8'b00001100;
        rContents[317] = 8'b00000000;
        rContents[318] = 8'b01100000;
        rContents[319] = 8'b00000100;
        rContents[320] = 8'b10000100;
        rContents[321] = 8'b00001010;
        rContents[322] = 8'b10000010;
        rContents[323] = 8'b10000000;
        rContents[324] = 8'b10000010;
        rContents[325] = 8'b10000000;
        rContents[326] = 8'b10000000;
        rContents[327] = 8'b10000000;
        rContents[328] = 8'b10000010;
        rContents[329] = 8'b00010000;
        rContents[330] = 8'b00000010;
        rContents[331] = 8'b10000100;
        rContents[332] = 8'b10000000;
        rContents[333] = 8'b10010010;
        rContents[334] = 8'b10000010;
        rContents[335] = 8'b10000010;
        rContents[336] = 8'b10000010;
        rContents[337] = 8'b10000010;
        rContents[338] = 8'b10000010;
        rContents[339] = 8'b10000000;
        rContents[340] = 8'b00010000;
        rContents[341] = 8'b10000010;
        rContents[342] = 8'b01000010;
        rContents[343] = 8'b10000010;
        rContents[344] = 8'b10000010;
        rContents[345] = 8'b10000010;
        rContents[346] = 8'b00000010;
        rContents[347] = 8'b00100000;
        rContents[348] = 8'b10000000;
        rContents[349] = 8'b00001000;
        rContents[350] = 8'b00101000;
        rContents[351] = 8'b00000000;
        rContents[352] = 8'b00010000;
        rContents[353] = 8'b00000000;
        rContents[354] = 8'b10000000;
        rContents[355] = 8'b00000000;
        rContents[356] = 8'b00000010;
        rContents[357] = 8'b00000000;
        rContents[358] = 8'b10000010;
        rContents[359] = 8'b00000000;
        rContents[360] = 8'b10000000;
        rContents[361] = 8'b00000000;
        rContents[362] = 8'b00000000;
        rContents[363] = 8'b10000000;
        rContents[364] = 8'b00010000;
        rContents[365] = 8'b00000000;
        rContents[366] = 8'b00000000;
        rContents[367] = 8'b00000000;
        rContents[368] = 8'b00000000;
        rContents[369] = 8'b00000000;
        rContents[370] = 8'b00000000;
        rContents[371] = 8'b00000000;
        rContents[372] = 8'b10000000;
        rContents[373] = 8'b00000000;
        rContents[374] = 8'b00000000;
        rContents[375] = 8'b00000000;
        rContents[376] = 8'b00000000;
        rContents[377] = 8'b00000000;
        rContents[378] = 8'b00000000;
        rContents[379] = 8'b00100000;
        rContents[380] = 8'b00010000;
        rContents[381] = 8'b00001000;
        rContents[382] = 8'b00000000;
        rContents[383] = 8'b00000000;
        rContents[384] = 8'b00000000;
        rContents[385] = 8'b11111111;
        rContents[386] = 8'b11111111;
        rContents[387] = 8'b11110000;
        rContents[388] = 8'b00001111;
        rContents[389] = 8'b11110000;
        rContents[390] = 8'b00001111;
        rContents[391] = 8'b00000000;
        rContents[392] = 8'b00000000;
        rContents[393] = 8'b11110000;
        rContents[394] = 8'b00001111;
        rContents[395] = 8'b11111111;
        rContents[396] = 8'b00000000;
        rContents[397] = 8'b00011000;
        rContents[398] = 8'b00000000;
        rContents[399] = 8'b00011000;
        rContents[400] = 8'b00011000;
        rContents[401] = 8'b00000000;
        rContents[402] = 8'b00000000;
        rContents[403] = 8'b00011000;
        rContents[404] = 8'b00000000;
        rContents[405] = 8'b00011000;
        rContents[406] = 8'b00011000;
        rContents[407] = 8'b00011000;
        rContents[408] = 8'b00100100;
        rContents[409] = 8'b00000000;
        rContents[410] = 8'b00100100;
        rContents[411] = 8'b00100100;
        rContents[412] = 8'b00000000;
        rContents[413] = 8'b00000000;
        rContents[414] = 8'b00100100;
        rContents[415] = 8'b00000000;
        rContents[416] = 8'b00100100;
        rContents[417] = 8'b00100100;
        rContents[418] = 8'b01000100;
        rContents[419] = 8'b00000000;
        rContents[420] = 8'b00000000;
        rContents[421] = 8'b10000010;
        rContents[422] = 8'b10000010;
        rContents[423] = 8'b00000100;
        rContents[424] = 8'b00000000;
        rContents[425] = 8'b00000000;
        rContents[426] = 8'b00000000;
        rContents[427] = 8'b00000000;
        rContents[428] = 8'b00000000;
        rContents[429] = 8'b00000000;
        rContents[430] = 8'b00000000;
        rContents[431] = 8'b00000000;
        rContents[432] = 8'b00000000;
        rContents[433] = 8'b00000000;
        rContents[434] = 8'b00000000;
        rContents[435] = 8'b00000000;
        rContents[436] = 8'b00000000;
        rContents[437] = 8'b00000000;
        rContents[438] = 8'b00000000;
        rContents[439] = 8'b00000000;
        rContents[440] = 8'b00000000;
        rContents[441] = 8'b00000000;
        rContents[442] = 8'b00000000;
        rContents[443] = 8'b00000000;
        rContents[444] = 8'b00000000;
        rContents[445] = 8'b00000000;
        rContents[446] = 8'b00000000;
        rContents[447] = 8'b00000000;
        rContents[448] = 8'b00000000;
        rContents[449] = 8'b00000000;
        rContents[450] = 8'b00000000;
        rContents[451] = 8'b00000000;
        rContents[452] = 8'b00000000;
        rContents[453] = 8'b00000000;
        rContents[454] = 8'b00000000;
        rContents[455] = 8'b00000000;
        rContents[456] = 8'b00000000;
        rContents[457] = 8'b00000000;
        rContents[458] = 8'b00000000;
        rContents[459] = 8'b00000000;
        rContents[460] = 8'b00000000;
        rContents[461] = 8'b00000000;
        rContents[462] = 8'b00000000;
        rContents[463] = 8'b00000000;
        rContents[464] = 8'b00000000;
        rContents[465] = 8'b00000000;
        rContents[466] = 8'b00000000;
        rContents[467] = 8'b00000000;
        rContents[468] = 8'b00000000;
        rContents[469] = 8'b00000000;
        rContents[470] = 8'b00000000;
        rContents[471] = 8'b00000000;
        rContents[472] = 8'b00000000;
        rContents[473] = 8'b00000000;
        rContents[474] = 8'b00000000;
        rContents[475] = 8'b00000000;
        rContents[476] = 8'b00000000;
        rContents[477] = 8'b00000000;
        rContents[478] = 8'b00000000;
        rContents[479] = 8'b00000000;
        rContents[480] = 8'b00000000;
        rContents[481] = 8'b00000000;
        rContents[482] = 8'b00000000;
        rContents[483] = 8'b00000000;
        rContents[484] = 8'b00000000;
        rContents[485] = 8'b00000000;
        rContents[486] = 8'b00000000;
        rContents[487] = 8'b00000000;
        rContents[488] = 8'b00000000;
        rContents[489] = 8'b00000000;
        rContents[490] = 8'b00000000;
        rContents[491] = 8'b00000000;
        rContents[492] = 8'b00000000;
        rContents[493] = 8'b00000000;
        rContents[494] = 8'b00000000;
        rContents[495] = 8'b00000000;
        rContents[496] = 8'b00000000;
        rContents[497] = 8'b00000000;
        rContents[498] = 8'b00000000;
        rContents[499] = 8'b00000000;
        rContents[500] = 8'b00000000;
        rContents[501] = 8'b00000000;
        rContents[502] = 8'b00000000;
        rContents[503] = 8'b00000000;
        rContents[504] = 8'b00000000;
        rContents[505] = 8'b00000000;
        rContents[506] = 8'b00000000;
        rContents[507] = 8'b00000000;
        rContents[508] = 8'b00000000;
        rContents[509] = 8'b00000000;
        rContents[510] = 8'b00000000;
        rContents[511] = 8'b00000000;
        rContents[512] = 8'b01010101;
        rContents[513] = 8'b10101010;
        rContents[514] = 8'b01010101;
        rContents[515] = 8'b11111111;
        rContents[516] = 8'b11111111;
        rContents[517] = 8'b00000000;
        rContents[518] = 8'b11111110;
        rContents[519] = 8'b10000010;
        rContents[520] = 8'b00010000;
        rContents[521] = 8'b10000010;
        rContents[522] = 8'b11111110;
        rContents[523] = 8'b11111110;
        rContents[524] = 8'b00111000;
        rContents[525] = 8'b00111000;
        rContents[526] = 8'b00111000;
        rContents[527] = 8'b10000010;
        rContents[528] = 8'b10010010;
        rContents[529] = 8'b11111110;
        rContents[530] = 8'b00100000;
        rContents[531] = 8'b00100010;
        rContents[532] = 8'b01111100;
        rContents[533] = 8'b00010000;
        rContents[534] = 8'b00100000;
        rContents[535] = 8'b00001000;
        rContents[536] = 8'b11111000;
        rContents[537] = 8'b00111110;
        rContents[538] = 8'b01111100;
        rContents[539] = 8'b10001010;
        rContents[540] = 8'b01111100;
        rContents[541] = 8'b00000000;
        rContents[542] = 8'b01111100;
        rContents[543] = 8'b01100000;
        rContents[544] = 8'b00000000;
        rContents[545] = 8'b00010000;
        rContents[546] = 8'b00000000;
        rContents[547] = 8'b11111110;
        rContents[548] = 8'b10010000;
        rContents[549] = 8'b11100100;
        rContents[550] = 8'b10000010;
        rContents[551] = 8'b00000000;
        rContents[552] = 8'b00100000;
        rContents[553] = 8'b00001000;
        rContents[554] = 8'b00010000;
        rContents[555] = 8'b00010000;
        rContents[556] = 8'b00000000;
        rContents[557] = 8'b00000000;
        rContents[558] = 8'b00000000;
        rContents[559] = 8'b00000100;
        rContents[560] = 8'b10000010;
        rContents[561] = 8'b00010000;
        rContents[562] = 8'b10000100;
        rContents[563] = 8'b00000010;
        rContents[564] = 8'b10000010;
        rContents[565] = 8'b10000000;
        rContents[566] = 8'b10000000;
        rContents[567] = 8'b00000010;
        rContents[568] = 8'b10000010;
        rContents[569] = 8'b10000010;
        rContents[570] = 8'b00000000;
        rContents[571] = 8'b00000000;
        rContents[572] = 8'b00010000;
        rContents[573] = 8'b00000000;
        rContents[574] = 8'b00010000;
        rContents[575] = 8'b00000100;
        rContents[576] = 8'b10111100;
        rContents[577] = 8'b00001010;
        rContents[578] = 8'b10000010;
        rContents[579] = 8'b10000000;
        rContents[580] = 8'b10000010;
        rContents[581] = 8'b10000000;
        rContents[582] = 8'b10000000;
        rContents[583] = 8'b10000000;
        rContents[584] = 8'b10000010;
        rContents[585] = 8'b00010000;
        rContents[586] = 8'b00000010;
        rContents[587] = 8'b10001000;
        rContents[588] = 8'b10000000;
        rContents[589] = 8'b10010010;
        rContents[590] = 8'b11000010;
        rContents[591] = 8'b10000010;
        rContents[592] = 8'b10000010;
        rContents[593] = 8'b10000010;
        rContents[594] = 8'b10000010;
        rContents[595] = 8'b10000000;
        rContents[596] = 8'b00010000;
        rContents[597] = 8'b10000010;
        rContents[598] = 8'b01000010;
        rContents[599] = 8'b10000010;
        rContents[600] = 8'b01000100;
        rContents[601] = 8'b01000100;
        rContents[602] = 8'b00000100;
        rContents[603] = 8'b00100000;
        rContents[604] = 8'b01000000;
        rContents[605] = 8'b00001000;
        rContents[606] = 8'b01000100;
        rContents[607] = 8'b00000000;
        rContents[608] = 8'b00000000;
        rContents[609] = 8'b00000000;
        rContents[610] = 8'b10000000;
        rContents[611] = 8'b00000000;
        rContents[612] = 8'b00000010;
        rContents[613] = 8'b00000000;
        rContents[614] = 8'b10000000;
        rContents[615] = 8'b00000000;
        rContents[616] = 8'b10000000;
        rContents[617] = 8'b00010000;
        rContents[618] = 8'b00001000;
        rContents[619] = 8'b10000000;
        rContents[620] = 8'b00010000;
        rContents[621] = 8'b00000000;
        rContents[622] = 8'b00000000;
        rContents[623] = 8'b00000000;
        rContents[624] = 8'b00000000;
        rContents[625] = 8'b00000000;
        rContents[626] = 8'b00000000;
        rContents[627] = 8'b00000000;
        rContents[628] = 8'b10000000;
        rContents[629] = 8'b00000000;
        rContents[630] = 8'b00000000;
        rContents[631] = 8'b00000000;
        rContents[632] = 8'b00000000;
        rContents[633] = 8'b00000000;
        rContents[634] = 8'b00000000;
        rContents[635] = 8'b00100000;
        rContents[636] = 8'b00010000;
        rContents[637] = 8'b00001000;
        rContents[638] = 8'b00000000;
        rContents[639] = 8'b00010000;
        rContents[640] = 8'b00010000;
        rContents[641] = 8'b11111111;
        rContents[642] = 8'b11111111;
        rContents[643] = 8'b11110000;
        rContents[644] = 8'b00001111;
        rContents[645] = 8'b11110000;
        rContents[646] = 8'b00001111;
        rContents[647] = 8'b00000000;
        rContents[648] = 8'b00000000;
        rContents[649] = 8'b11110000;
        rContents[650] = 8'b00001111;
        rContents[651] = 8'b11111111;
        rContents[652] = 8'b00000000;
        rContents[653] = 8'b00011000;
        rContents[654] = 8'b00000000;
        rContents[655] = 8'b00011000;
        rContents[656] = 8'b00011000;
        rContents[657] = 8'b00000000;
        rContents[658] = 8'b00000000;
        rContents[659] = 8'b00011000;
        rContents[660] = 8'b00000000;
        rContents[661] = 8'b00011000;
        rContents[662] = 8'b00011000;
        rContents[663] = 8'b00011000;
        rContents[664] = 8'b00100100;
        rContents[665] = 8'b00000000;
        rContents[666] = 8'b00100100;
        rContents[667] = 8'b00100100;
        rContents[668] = 8'b00000000;
        rContents[669] = 8'b00000000;
        rContents[670] = 8'b00100100;
        rContents[671] = 8'b00000000;
        rContents[672] = 8'b00100100;
        rContents[673] = 8'b00100100;
        rContents[674] = 8'b10000010;
        rContents[675] = 8'b00000000;
        rContents[676] = 8'b00000000;
        rContents[677] = 8'b10000010;
        rContents[678] = 8'b01000000;
        rContents[679] = 8'b00000100;
        rContents[680] = 8'b00000000;
        rContents[681] = 8'b00000000;
        rContents[682] = 8'b00000000;
        rContents[683] = 8'b00000000;
        rContents[684] = 8'b00000000;
        rContents[685] = 8'b00000000;
        rContents[686] = 8'b00000000;
        rContents[687] = 8'b00000000;
        rContents[688] = 8'b00000000;
        rContents[689] = 8'b00000000;
        rContents[690] = 8'b00000000;
        rContents[691] = 8'b00000000;
        rContents[692] = 8'b00000000;
        rContents[693] = 8'b00000000;
        rContents[694] = 8'b00000000;
        rContents[695] = 8'b00000000;
        rContents[696] = 8'b00000000;
        rContents[697] = 8'b00000000;
        rContents[698] = 8'b00000000;
        rContents[699] = 8'b00000000;
        rContents[700] = 8'b00000000;
        rContents[701] = 8'b00000000;
        rContents[702] = 8'b00000000;
        rContents[703] = 8'b00000000;
        rContents[704] = 8'b00000000;
        rContents[705] = 8'b00000000;
        rContents[706] = 8'b00000000;
        rContents[707] = 8'b00000000;
        rContents[708] = 8'b00000000;
        rContents[709] = 8'b00000000;
        rContents[710] = 8'b00000000;
        rContents[711] = 8'b00000000;
        rContents[712] = 8'b00000000;
        rContents[713] = 8'b00000000;
        rContents[714] = 8'b00000000;
        rContents[715] = 8'b00000000;
        rContents[716] = 8'b00000000;
        rContents[717] = 8'b00000000;
        rContents[718] = 8'b00000000;
        rContents[719] = 8'b00000000;
        rContents[720] = 8'b00000000;
        rContents[721] = 8'b00000000;
        rContents[722] = 8'b00000000;
        rContents[723] = 8'b00000000;
        rContents[724] = 8'b00000000;
        rContents[725] = 8'b00000000;
        rContents[726] = 8'b00000000;
        rContents[727] = 8'b00000000;
        rContents[728] = 8'b00000000;
        rContents[729] = 8'b00000000;
        rContents[730] = 8'b00000000;
        rContents[731] = 8'b00000000;
        rContents[732] = 8'b00000000;
        rContents[733] = 8'b00000000;
        rContents[734] = 8'b00000000;
        rContents[735] = 8'b00000000;
        rContents[736] = 8'b00000000;
        rContents[737] = 8'b00000000;
        rContents[738] = 8'b00000000;
        rContents[739] = 8'b00000000;
        rContents[740] = 8'b00000000;
        rContents[741] = 8'b00000000;
        rContents[742] = 8'b00000000;
        rContents[743] = 8'b00000000;
        rContents[744] = 8'b00000000;
        rContents[745] = 8'b00000000;
        rContents[746] = 8'b00000000;
        rContents[747] = 8'b00000000;
        rContents[748] = 8'b00000000;
        rContents[749] = 8'b00000000;
        rContents[750] = 8'b00000000;
        rContents[751] = 8'b00000000;
        rContents[752] = 8'b00000000;
        rContents[753] = 8'b00000000;
        rContents[754] = 8'b00000000;
        rContents[755] = 8'b00000000;
        rContents[756] = 8'b00000000;
        rContents[757] = 8'b00000000;
        rContents[758] = 8'b00000000;
        rContents[759] = 8'b00000000;
        rContents[760] = 8'b00000000;
        rContents[761] = 8'b00000000;
        rContents[762] = 8'b00000000;
        rContents[763] = 8'b00000000;
        rContents[764] = 8'b00000000;
        rContents[765] = 8'b00000000;
        rContents[766] = 8'b00000000;
        rContents[767] = 8'b00000000;
        rContents[768] = 8'b01010101;
        rContents[769] = 8'b10101010;
        rContents[770] = 8'b11111111;
        rContents[771] = 8'b10101010;
        rContents[772] = 8'b11111111;
        rContents[773] = 8'b00000000;
        rContents[774] = 8'b11111110;
        rContents[775] = 8'b10000010;
        rContents[776] = 8'b00010000;
        rContents[777] = 8'b10101010;
        rContents[778] = 8'b11010110;
        rContents[779] = 8'b11111110;
        rContents[780] = 8'b01111100;
        rContents[781] = 8'b11111110;
        rContents[782] = 8'b01111100;
        rContents[783] = 8'b10010010;
        rContents[784] = 8'b10101010;
        rContents[785] = 8'b11101110;
        rContents[786] = 8'b00100000;
        rContents[787] = 8'b00100010;
        rContents[788] = 8'b00010000;
        rContents[789] = 8'b00010000;
        rContents[790] = 8'b01100000;
        rContents[791] = 8'b00001100;
        rContents[792] = 8'b11111100;
        rContents[793] = 8'b01111110;
        rContents[794] = 8'b00010000;
        rContents[795] = 8'b10001010;
        rContents[796] = 8'b01111100;
        rContents[797] = 8'b11111110;
        rContents[798] = 8'b00010000;
        rContents[799] = 8'b00111000;
        rContents[800] = 8'b00000000;
        rContents[801] = 8'b00010000;
        rContents[802] = 8'b00000000;
        rContents[803] = 8'b01000100;
        rContents[804] = 8'b10010000;
        rContents[805] = 8'b00001000;
        rContents[806] = 8'b10000010;
        rContents[807] = 8'b00000000;
        rContents[808] = 8'b00100000;
        rContents[809] = 8'b00001000;
        rContents[810] = 8'b00000000;
        rContents[811] = 8'b00010000;
        rContents[812] = 8'b00000000;
        rContents[813] = 8'b00000000;
        rContents[814] = 8'b00000000;
        rContents[815] = 8'b00001000;
        rContents[816] = 8'b10010010;
        rContents[817] = 8'b00010000;
        rContents[818] = 8'b00001000;
        rContents[819] = 8'b00000010;
        rContents[820] = 8'b10000010;
        rContents[821] = 8'b10000000;
        rContents[822] = 8'b10000000;
        rContents[823] = 8'b00000100;
        rContents[824] = 8'b10000010;
        rContents[825] = 8'b10000010;
        rContents[826] = 8'b00000000;
        rContents[827] = 8'b00000000;
        rContents[828] = 8'b01100000;
        rContents[829] = 8'b11111110;
        rContents[830] = 8'b00001100;
        rContents[831] = 8'b00000100;
        rContents[832] = 8'b10100100;
        rContents[833] = 8'b00010010;
        rContents[834] = 8'b10000010;
        rContents[835] = 8'b10000000;
        rContents[836] = 8'b10000010;
        rContents[837] = 8'b10000000;
        rContents[838] = 8'b10000000;
        rContents[839] = 8'b10000000;
        rContents[840] = 8'b10000010;
        rContents[841] = 8'b00010000;
        rContents[842] = 8'b00000010;
        rContents[843] = 8'b10010000;
        rContents[844] = 8'b10000000;
        rContents[845] = 8'b10010010;
        rContents[846] = 8'b10100010;
        rContents[847] = 8'b10000010;
        rContents[848] = 8'b10000010;
        rContents[849] = 8'b10000010;
        rContents[850] = 8'b10000010;
        rContents[851] = 8'b10000000;
        rContents[852] = 8'b00010000;
        rContents[853] = 8'b10000010;
        rContents[854] = 8'b00100010;
        rContents[855] = 8'b10000010;
        rContents[856] = 8'b00101000;
        rContents[857] = 8'b00101000;
        rContents[858] = 8'b00001000;
        rContents[859] = 8'b00100000;
        rContents[860] = 8'b00100000;
        rContents[861] = 8'b00001000;
        rContents[862] = 8'b00000000;
        rContents[863] = 8'b00000000;
        rContents[864] = 8'b00000000;
        rContents[865] = 8'b00000000;
        rContents[866] = 8'b10000000;
        rContents[867] = 8'b00000000;
        rContents[868] = 8'b00000010;
        rContents[869] = 8'b00000000;
        rContents[870] = 8'b10000000;
        rContents[871] = 8'b00000000;
        rContents[872] = 8'b10000000;
        rContents[873] = 8'b00000000;
        rContents[874] = 8'b00000000;
        rContents[875] = 8'b10000000;
        rContents[876] = 8'b00010000;
        rContents[877] = 8'b00000000;
        rContents[878] = 8'b00000000;
        rContents[879] = 8'b00000000;
        rContents[880] = 8'b00000000;
        rContents[881] = 8'b00000000;
        rContents[882] = 8'b00000000;
        rContents[883] = 8'b00000000;
        rContents[884] = 8'b10000000;
        rContents[885] = 8'b00000000;
        rContents[886] = 8'b00000000;
        rContents[887] = 8'b00000000;
        rContents[888] = 8'b00000000;
        rContents[889] = 8'b00000000;
        rContents[890] = 8'b00000000;
        rContents[891] = 8'b00100000;
        rContents[892] = 8'b00010000;
        rContents[893] = 8'b00001000;
        rContents[894] = 8'b01100000;
        rContents[895] = 8'b00010000;
        rContents[896] = 8'b00010000;
        rContents[897] = 8'b11111111;
        rContents[898] = 8'b11111111;
        rContents[899] = 8'b11110000;
        rContents[900] = 8'b00001111;
        rContents[901] = 8'b11110000;
        rContents[902] = 8'b00001111;
        rContents[903] = 8'b00000000;
        rContents[904] = 8'b00000000;
        rContents[905] = 8'b11110000;
        rContents[906] = 8'b00001111;
        rContents[907] = 8'b11111111;
        rContents[908] = 8'b00000000;
        rContents[909] = 8'b00011000;
        rContents[910] = 8'b00000000;
        rContents[911] = 8'b00011000;
        rContents[912] = 8'b00011000;
        rContents[913] = 8'b00000000;
        rContents[914] = 8'b00000000;
        rContents[915] = 8'b00011000;
        rContents[916] = 8'b00000000;
        rContents[917] = 8'b00011000;
        rContents[918] = 8'b00011000;
        rContents[919] = 8'b00011000;
        rContents[920] = 8'b00100100;
        rContents[921] = 8'b00000000;
        rContents[922] = 8'b00100100;
        rContents[923] = 8'b00100100;
        rContents[924] = 8'b00000000;
        rContents[925] = 8'b00000000;
        rContents[926] = 8'b00100100;
        rContents[927] = 8'b00000000;
        rContents[928] = 8'b00100100;
        rContents[929] = 8'b00100100;
        rContents[930] = 8'b10000010;
        rContents[931] = 8'b00000000;
        rContents[932] = 8'b00000000;
        rContents[933] = 8'b11111100;
        rContents[934] = 8'b00100000;
        rContents[935] = 8'b00000100;
        rContents[936] = 8'b00000000;
        rContents[937] = 8'b00000000;
        rContents[938] = 8'b00000000;
        rContents[939] = 8'b00000000;
        rContents[940] = 8'b00000000;
        rContents[941] = 8'b00000000;
        rContents[942] = 8'b00000000;
        rContents[943] = 8'b00000000;
        rContents[944] = 8'b00000000;
        rContents[945] = 8'b00000000;
        rContents[946] = 8'b00000000;
        rContents[947] = 8'b00000000;
        rContents[948] = 8'b00000000;
        rContents[949] = 8'b00000000;
        rContents[950] = 8'b00000000;
        rContents[951] = 8'b00000000;
        rContents[952] = 8'b00000000;
        rContents[953] = 8'b00000000;
        rContents[954] = 8'b00000000;
        rContents[955] = 8'b00000000;
        rContents[956] = 8'b00000000;
        rContents[957] = 8'b00000000;
        rContents[958] = 8'b00000000;
        rContents[959] = 8'b00000000;
        rContents[960] = 8'b00000000;
        rContents[961] = 8'b00000000;
        rContents[962] = 8'b00000000;
        rContents[963] = 8'b00000000;
        rContents[964] = 8'b00000000;
        rContents[965] = 8'b00000000;
        rContents[966] = 8'b00000000;
        rContents[967] = 8'b00000000;
        rContents[968] = 8'b00000000;
        rContents[969] = 8'b00000000;
        rContents[970] = 8'b00000000;
        rContents[971] = 8'b00000000;
        rContents[972] = 8'b00000000;
        rContents[973] = 8'b00000000;
        rContents[974] = 8'b00000000;
        rContents[975] = 8'b00000000;
        rContents[976] = 8'b00000000;
        rContents[977] = 8'b00000000;
        rContents[978] = 8'b00000000;
        rContents[979] = 8'b00000000;
        rContents[980] = 8'b00000000;
        rContents[981] = 8'b00000000;
        rContents[982] = 8'b00000000;
        rContents[983] = 8'b00000000;
        rContents[984] = 8'b00000000;
        rContents[985] = 8'b00000000;
        rContents[986] = 8'b00000000;
        rContents[987] = 8'b00000000;
        rContents[988] = 8'b00000000;
        rContents[989] = 8'b00000000;
        rContents[990] = 8'b00000000;
        rContents[991] = 8'b00000000;
        rContents[992] = 8'b00000000;
        rContents[993] = 8'b00000000;
        rContents[994] = 8'b00000000;
        rContents[995] = 8'b00000000;
        rContents[996] = 8'b00000000;
        rContents[997] = 8'b00000000;
        rContents[998] = 8'b00000000;
        rContents[999] = 8'b00000000;
        rContents[1000] = 8'b00000000;
        rContents[1001] = 8'b00000000;
        rContents[1002] = 8'b00000000;
        rContents[1003] = 8'b00000000;
        rContents[1004] = 8'b00000000;
        rContents[1005] = 8'b00000000;
        rContents[1006] = 8'b00000000;
        rContents[1007] = 8'b00000000;
        rContents[1008] = 8'b00000000;
        rContents[1009] = 8'b00000000;
        rContents[1010] = 8'b00000000;
        rContents[1011] = 8'b00000000;
        rContents[1012] = 8'b00000000;
        rContents[1013] = 8'b00000000;
        rContents[1014] = 8'b00000000;
        rContents[1015] = 8'b00000000;
        rContents[1016] = 8'b00000000;
        rContents[1017] = 8'b00000000;
        rContents[1018] = 8'b00000000;
        rContents[1019] = 8'b00000000;
        rContents[1020] = 8'b00000000;
        rContents[1021] = 8'b00000000;
        rContents[1022] = 8'b00000000;
        rContents[1023] = 8'b00000000;
        rContents[1024] = 8'b01010101;
        rContents[1025] = 8'b10101010;
        rContents[1026] = 8'b01010101;
        rContents[1027] = 8'b11111111;
        rContents[1028] = 8'b11111111;
        rContents[1029] = 8'b00000000;
        rContents[1030] = 8'b11111110;
        rContents[1031] = 8'b10000010;
        rContents[1032] = 8'b00010000;
        rContents[1033] = 8'b10000010;
        rContents[1034] = 8'b11111110;
        rContents[1035] = 8'b01111100;
        rContents[1036] = 8'b11111110;
        rContents[1037] = 8'b11111110;
        rContents[1038] = 8'b11111110;
        rContents[1039] = 8'b10111010;
        rContents[1040] = 8'b11000110;
        rContents[1041] = 8'b11000110;
        rContents[1042] = 8'b00100000;
        rContents[1043] = 8'b00100010;
        rContents[1044] = 8'b00010000;
        rContents[1045] = 8'b00010000;
        rContents[1046] = 8'b11111110;
        rContents[1047] = 8'b11111110;
        rContents[1048] = 8'b11111110;
        rContents[1049] = 8'b11111110;
        rContents[1050] = 8'b00010000;
        rContents[1051] = 8'b11111110;
        rContents[1052] = 8'b11111110;
        rContents[1053] = 8'b11111110;
        rContents[1054] = 8'b00010000;
        rContents[1055] = 8'b00101000;
        rContents[1056] = 8'b00000000;
        rContents[1057] = 8'b00010000;
        rContents[1058] = 8'b00000000;
        rContents[1059] = 8'b01000100;
        rContents[1060] = 8'b11111110;
        rContents[1061] = 8'b00010000;
        rContents[1062] = 8'b01101100;
        rContents[1063] = 8'b00000000;
        rContents[1064] = 8'b00100000;
        rContents[1065] = 8'b00001000;
        rContents[1066] = 8'b00000000;
        rContents[1067] = 8'b00010000;
        rContents[1068] = 8'b00000000;
        rContents[1069] = 8'b00000000;
        rContents[1070] = 8'b00000000;
        rContents[1071] = 8'b00010000;
        rContents[1072] = 8'b10010010;
        rContents[1073] = 8'b00010000;
        rContents[1074] = 8'b00010000;
        rContents[1075] = 8'b00011110;
        rContents[1076] = 8'b11111110;
        rContents[1077] = 8'b11111100;
        rContents[1078] = 8'b11111100;
        rContents[1079] = 8'b00000100;
        rContents[1080] = 8'b01111100;
        rContents[1081] = 8'b01111110;
        rContents[1082] = 8'b00000000;
        rContents[1083] = 8'b00000000;
        rContents[1084] = 8'b10000000;
        rContents[1085] = 8'b00000000;
        rContents[1086] = 8'b00000010;
        rContents[1087] = 8'b00011100;
        rContents[1088] = 8'b10100100;
        rContents[1089] = 8'b00111110;
        rContents[1090] = 8'b11111100;
        rContents[1091] = 8'b10000000;
        rContents[1092] = 8'b10000010;
        rContents[1093] = 8'b11111110;
        rContents[1094] = 8'b11111110;
        rContents[1095] = 8'b10001110;
        rContents[1096] = 8'b11111110;
        rContents[1097] = 8'b00010000;
        rContents[1098] = 8'b00000010;
        rContents[1099] = 8'b11100000;
        rContents[1100] = 8'b10000000;
        rContents[1101] = 8'b10010010;
        rContents[1102] = 8'b10010010;
        rContents[1103] = 8'b10000010;
        rContents[1104] = 8'b11111110;
        rContents[1105] = 8'b10000010;
        rContents[1106] = 8'b11111110;
        rContents[1107] = 8'b11111110;
        rContents[1108] = 8'b00010000;
        rContents[1109] = 8'b10000010;
        rContents[1110] = 8'b00100010;
        rContents[1111] = 8'b10010010;
        rContents[1112] = 8'b00010000;
        rContents[1113] = 8'b00010000;
        rContents[1114] = 8'b00010000;
        rContents[1115] = 8'b00100000;
        rContents[1116] = 8'b00010000;
        rContents[1117] = 8'b00001000;
        rContents[1118] = 8'b00000000;
        rContents[1119] = 8'b00000000;
        rContents[1120] = 8'b00000000;
        rContents[1121] = 8'b11111110;
        rContents[1122] = 8'b11111110;
        rContents[1123] = 8'b11111110;
        rContents[1124] = 8'b11111110;
        rContents[1125] = 8'b11111110;
        rContents[1126] = 8'b11110000;
        rContents[1127] = 8'b11111110;
        rContents[1128] = 8'b11111110;
        rContents[1129] = 8'b00010000;
        rContents[1130] = 8'b00001000;
        rContents[1131] = 8'b10000110;
        rContents[1132] = 8'b00010000;
        rContents[1133] = 8'b11111110;
        rContents[1134] = 8'b11111110;
        rContents[1135] = 8'b11111110;
        rContents[1136] = 8'b11111110;
        rContents[1137] = 8'b11111110;
        rContents[1138] = 8'b11111110;
        rContents[1139] = 8'b11111110;
        rContents[1140] = 8'b11111110;
        rContents[1141] = 8'b10000010;
        rContents[1142] = 8'b10000010;
        rContents[1143] = 8'b10000010;
        rContents[1144] = 8'b11000110;
        rContents[1145] = 8'b10000010;
        rContents[1146] = 8'b11111110;
        rContents[1147] = 8'b01000000;
        rContents[1148] = 8'b00010000;
        rContents[1149] = 8'b00000100;
        rContents[1150] = 8'b10010010;
        rContents[1151] = 8'b00010000;
        rContents[1152] = 8'b00011100;
        rContents[1153] = 8'b11111111;
        rContents[1154] = 8'b11111111;
        rContents[1155] = 8'b11110000;
        rContents[1156] = 8'b00001111;
        rContents[1157] = 8'b11110000;
        rContents[1158] = 8'b00001111;
        rContents[1159] = 8'b00000000;
        rContents[1160] = 8'b00000000;
        rContents[1161] = 8'b11110000;
        rContents[1162] = 8'b00001111;
        rContents[1163] = 8'b11111111;
        rContents[1164] = 8'b00000000;
        rContents[1165] = 8'b00011000;
        rContents[1166] = 8'b00000000;
        rContents[1167] = 8'b00011000;
        rContents[1168] = 8'b00011000;
        rContents[1169] = 8'b00000000;
        rContents[1170] = 8'b00000000;
        rContents[1171] = 8'b00011000;
        rContents[1172] = 8'b00000000;
        rContents[1173] = 8'b00011000;
        rContents[1174] = 8'b00011000;
        rContents[1175] = 8'b00011000;
        rContents[1176] = 8'b00100100;
        rContents[1177] = 8'b11111111;
        rContents[1178] = 8'b11100111;
        rContents[1179] = 8'b11100111;
        rContents[1180] = 8'b11111111;
        rContents[1181] = 8'b11111100;
        rContents[1182] = 8'b11100100;
        rContents[1183] = 8'b00111111;
        rContents[1184] = 8'b11100100;
        rContents[1185] = 8'b00100111;
        rContents[1186] = 8'b10000010;
        rContents[1187] = 8'b11111110;
        rContents[1188] = 8'b01110010;
        rContents[1189] = 8'b10000010;
        rContents[1190] = 8'b00010000;
        rContents[1191] = 8'b11000100;
        rContents[1192] = 8'b00000000;
        rContents[1193] = 8'b00000000;
        rContents[1194] = 8'b00000000;
        rContents[1195] = 8'b00000000;
        rContents[1196] = 8'b00000000;
        rContents[1197] = 8'b00000000;
        rContents[1198] = 8'b00000000;
        rContents[1199] = 8'b00000000;
        rContents[1200] = 8'b00000000;
        rContents[1201] = 8'b00000000;
        rContents[1202] = 8'b00000000;
        rContents[1203] = 8'b00000000;
        rContents[1204] = 8'b00000000;
        rContents[1205] = 8'b00000000;
        rContents[1206] = 8'b00000000;
        rContents[1207] = 8'b00000000;
        rContents[1208] = 8'b00000000;
        rContents[1209] = 8'b00000000;
        rContents[1210] = 8'b00000000;
        rContents[1211] = 8'b00000000;
        rContents[1212] = 8'b00000000;
        rContents[1213] = 8'b00000000;
        rContents[1214] = 8'b00000000;
        rContents[1215] = 8'b00000000;
        rContents[1216] = 8'b00000000;
        rContents[1217] = 8'b00000000;
        rContents[1218] = 8'b00000000;
        rContents[1219] = 8'b00000000;
        rContents[1220] = 8'b00000000;
        rContents[1221] = 8'b00000000;
        rContents[1222] = 8'b00000000;
        rContents[1223] = 8'b00000000;
        rContents[1224] = 8'b00000000;
        rContents[1225] = 8'b00000000;
        rContents[1226] = 8'b00000000;
        rContents[1227] = 8'b00000000;
        rContents[1228] = 8'b00000000;
        rContents[1229] = 8'b00000000;
        rContents[1230] = 8'b00000000;
        rContents[1231] = 8'b00000000;
        rContents[1232] = 8'b00000000;
        rContents[1233] = 8'b00000000;
        rContents[1234] = 8'b00000000;
        rContents[1235] = 8'b00000000;
        rContents[1236] = 8'b00000000;
        rContents[1237] = 8'b00000000;
        rContents[1238] = 8'b00000000;
        rContents[1239] = 8'b00000000;
        rContents[1240] = 8'b00000000;
        rContents[1241] = 8'b00000000;
        rContents[1242] = 8'b00000000;
        rContents[1243] = 8'b00000000;
        rContents[1244] = 8'b00000000;
        rContents[1245] = 8'b00000000;
        rContents[1246] = 8'b00000000;
        rContents[1247] = 8'b00000000;
        rContents[1248] = 8'b00000000;
        rContents[1249] = 8'b00000000;
        rContents[1250] = 8'b00000000;
        rContents[1251] = 8'b00000000;
        rContents[1252] = 8'b00000000;
        rContents[1253] = 8'b00000000;
        rContents[1254] = 8'b00000000;
        rContents[1255] = 8'b00000000;
        rContents[1256] = 8'b00000000;
        rContents[1257] = 8'b00000000;
        rContents[1258] = 8'b00000000;
        rContents[1259] = 8'b00000000;
        rContents[1260] = 8'b00000000;
        rContents[1261] = 8'b00000000;
        rContents[1262] = 8'b00000000;
        rContents[1263] = 8'b00000000;
        rContents[1264] = 8'b00000000;
        rContents[1265] = 8'b00000000;
        rContents[1266] = 8'b00000000;
        rContents[1267] = 8'b00000000;
        rContents[1268] = 8'b00000000;
        rContents[1269] = 8'b00000000;
        rContents[1270] = 8'b00000000;
        rContents[1271] = 8'b00000000;
        rContents[1272] = 8'b00000000;
        rContents[1273] = 8'b00000000;
        rContents[1274] = 8'b00000000;
        rContents[1275] = 8'b00000000;
        rContents[1276] = 8'b00000000;
        rContents[1277] = 8'b00000000;
        rContents[1278] = 8'b00000000;
        rContents[1279] = 8'b00000000;
        rContents[1280] = 8'b01010101;
        rContents[1281] = 8'b10101010;
        rContents[1282] = 8'b11111111;
        rContents[1283] = 8'b10101010;
        rContents[1284] = 8'b11111111;
        rContents[1285] = 8'b00000000;
        rContents[1286] = 8'b11111110;
        rContents[1287] = 8'b10000010;
        rContents[1288] = 8'b00010000;
        rContents[1289] = 8'b10111010;
        rContents[1290] = 8'b11000110;
        rContents[1291] = 8'b01111100;
        rContents[1292] = 8'b01111100;
        rContents[1293] = 8'b11111110;
        rContents[1294] = 8'b01111100;
        rContents[1295] = 8'b10010010;
        rContents[1296] = 8'b10101010;
        rContents[1297] = 8'b11101110;
        rContents[1298] = 8'b01100000;
        rContents[1299] = 8'b01100110;
        rContents[1300] = 8'b00010000;
        rContents[1301] = 8'b00010000;
        rContents[1302] = 8'b01100000;
        rContents[1303] = 8'b00001100;
        rContents[1304] = 8'b11111100;
        rContents[1305] = 8'b01111110;
        rContents[1306] = 8'b00010000;
        rContents[1307] = 8'b00001010;
        rContents[1308] = 8'b11111110;
        rContents[1309] = 8'b01111100;
        rContents[1310] = 8'b01111100;
        rContents[1311] = 8'b00111000;
        rContents[1312] = 8'b00000000;
        rContents[1313] = 8'b00010000;
        rContents[1314] = 8'b00000000;
        rContents[1315] = 8'b01000100;
        rContents[1316] = 8'b00010010;
        rContents[1317] = 8'b00100000;
        rContents[1318] = 8'b00010000;
        rContents[1319] = 8'b00000000;
        rContents[1320] = 8'b00100000;
        rContents[1321] = 8'b00001000;
        rContents[1322] = 8'b00000000;
        rContents[1323] = 8'b11111110;
        rContents[1324] = 8'b00000000;
        rContents[1325] = 8'b11111110;
        rContents[1326] = 8'b00000000;
        rContents[1327] = 8'b00100000;
        rContents[1328] = 8'b10010010;
        rContents[1329] = 8'b00010000;
        rContents[1330] = 8'b00100000;
        rContents[1331] = 8'b00000010;
        rContents[1332] = 8'b00000010;
        rContents[1333] = 8'b00000010;
        rContents[1334] = 8'b10000010;
        rContents[1335] = 8'b00001000;
        rContents[1336] = 8'b10000010;
        rContents[1337] = 8'b00000010;
        rContents[1338] = 8'b00000000;
        rContents[1339] = 8'b00000000;
        rContents[1340] = 8'b01100000;
        rContents[1341] = 8'b00000000;
        rContents[1342] = 8'b00001100;
        rContents[1343] = 8'b00010000;
        rContents[1344] = 8'b10100100;
        rContents[1345] = 8'b00100010;
        rContents[1346] = 8'b10000010;
        rContents[1347] = 8'b10000000;
        rContents[1348] = 8'b10000010;
        rContents[1349] = 8'b10000000;
        rContents[1350] = 8'b10000000;
        rContents[1351] = 8'b10000010;
        rContents[1352] = 8'b10000010;
        rContents[1353] = 8'b00010000;
        rContents[1354] = 8'b00000010;
        rContents[1355] = 8'b10010000;
        rContents[1356] = 8'b10000000;
        rContents[1357] = 8'b10000010;
        rContents[1358] = 8'b10001010;
        rContents[1359] = 8'b10000010;
        rContents[1360] = 8'b10000000;
        rContents[1361] = 8'b10010010;
        rContents[1362] = 8'b11000000;
        rContents[1363] = 8'b00000010;
        rContents[1364] = 8'b00010000;
        rContents[1365] = 8'b10000010;
        rContents[1366] = 8'b00010010;
        rContents[1367] = 8'b10010010;
        rContents[1368] = 8'b00101000;
        rContents[1369] = 8'b00010000;
        rContents[1370] = 8'b00100000;
        rContents[1371] = 8'b00100000;
        rContents[1372] = 8'b00001000;
        rContents[1373] = 8'b00001000;
        rContents[1374] = 8'b00000000;
        rContents[1375] = 8'b00000000;
        rContents[1376] = 8'b00000000;
        rContents[1377] = 8'b00000010;
        rContents[1378] = 8'b10000010;
        rContents[1379] = 8'b10000000;
        rContents[1380] = 8'b10000010;
        rContents[1381] = 8'b10000010;
        rContents[1382] = 8'b10000000;
        rContents[1383] = 8'b10000010;
        rContents[1384] = 8'b10000010;
        rContents[1385] = 8'b00010000;
        rContents[1386] = 8'b00001000;
        rContents[1387] = 8'b10011000;
        rContents[1388] = 8'b00010000;
        rContents[1389] = 8'b10010010;
        rContents[1390] = 8'b10000010;
        rContents[1391] = 8'b10000010;
        rContents[1392] = 8'b10000010;
        rContents[1393] = 8'b10000010;
        rContents[1394] = 8'b10000000;
        rContents[1395] = 8'b10000000;
        rContents[1396] = 8'b10000000;
        rContents[1397] = 8'b10000010;
        rContents[1398] = 8'b01000010;
        rContents[1399] = 8'b10000010;
        rContents[1400] = 8'b00101000;
        rContents[1401] = 8'b10000010;
        rContents[1402] = 8'b00000100;
        rContents[1403] = 8'b00100000;
        rContents[1404] = 8'b00010000;
        rContents[1405] = 8'b00001000;
        rContents[1406] = 8'b00001100;
        rContents[1407] = 8'b00010000;
        rContents[1408] = 8'b00000100;
        rContents[1409] = 8'b11111111;
        rContents[1410] = 8'b11111111;
        rContents[1411] = 8'b11110000;
        rContents[1412] = 8'b00001111;
        rContents[1413] = 8'b11110000;
        rContents[1414] = 8'b00001111;
        rContents[1415] = 8'b00000000;
        rContents[1416] = 8'b00000000;
        rContents[1417] = 8'b11110000;
        rContents[1418] = 8'b00001111;
        rContents[1419] = 8'b11111111;
        rContents[1420] = 8'b00000000;
        rContents[1421] = 8'b00011000;
        rContents[1422] = 8'b11111111;
        rContents[1423] = 8'b11111111;
        rContents[1424] = 8'b11111111;
        rContents[1425] = 8'b11111111;
        rContents[1426] = 8'b11111000;
        rContents[1427] = 8'b11111000;
        rContents[1428] = 8'b00011111;
        rContents[1429] = 8'b00011111;
        rContents[1430] = 8'b11111000;
        rContents[1431] = 8'b00011111;
        rContents[1432] = 8'b00100100;
        rContents[1433] = 8'b00000000;
        rContents[1434] = 8'b00000000;
        rContents[1435] = 8'b00000000;
        rContents[1436] = 8'b00000000;
        rContents[1437] = 8'b00000100;
        rContents[1438] = 8'b00000100;
        rContents[1439] = 8'b00100000;
        rContents[1440] = 8'b00000100;
        rContents[1441] = 8'b00100000;
        rContents[1442] = 8'b10000010;
        rContents[1443] = 8'b01000100;
        rContents[1444] = 8'b10001100;
        rContents[1445] = 8'b10000010;
        rContents[1446] = 8'b00100000;
        rContents[1447] = 8'b00100100;
        rContents[1448] = 8'b00000000;
        rContents[1449] = 8'b00000000;
        rContents[1450] = 8'b00000000;
        rContents[1451] = 8'b00000000;
        rContents[1452] = 8'b00000000;
        rContents[1453] = 8'b00000000;
        rContents[1454] = 8'b00000000;
        rContents[1455] = 8'b00000000;
        rContents[1456] = 8'b00000000;
        rContents[1457] = 8'b00000000;
        rContents[1458] = 8'b00000000;
        rContents[1459] = 8'b00000000;
        rContents[1460] = 8'b00000000;
        rContents[1461] = 8'b00000000;
        rContents[1462] = 8'b00000000;
        rContents[1463] = 8'b00000000;
        rContents[1464] = 8'b00000000;
        rContents[1465] = 8'b00000000;
        rContents[1466] = 8'b00000000;
        rContents[1467] = 8'b00000000;
        rContents[1468] = 8'b00000000;
        rContents[1469] = 8'b00000000;
        rContents[1470] = 8'b00000000;
        rContents[1471] = 8'b00000000;
        rContents[1472] = 8'b00000000;
        rContents[1473] = 8'b00000000;
        rContents[1474] = 8'b00000000;
        rContents[1475] = 8'b00000000;
        rContents[1476] = 8'b00000000;
        rContents[1477] = 8'b00000000;
        rContents[1478] = 8'b00000000;
        rContents[1479] = 8'b00000000;
        rContents[1480] = 8'b00000000;
        rContents[1481] = 8'b00000000;
        rContents[1482] = 8'b00000000;
        rContents[1483] = 8'b00000000;
        rContents[1484] = 8'b00000000;
        rContents[1485] = 8'b00000000;
        rContents[1486] = 8'b00000000;
        rContents[1487] = 8'b00000000;
        rContents[1488] = 8'b00000000;
        rContents[1489] = 8'b00000000;
        rContents[1490] = 8'b00000000;
        rContents[1491] = 8'b00000000;
        rContents[1492] = 8'b00000000;
        rContents[1493] = 8'b00000000;
        rContents[1494] = 8'b00000000;
        rContents[1495] = 8'b00000000;
        rContents[1496] = 8'b00000000;
        rContents[1497] = 8'b00000000;
        rContents[1498] = 8'b00000000;
        rContents[1499] = 8'b00000000;
        rContents[1500] = 8'b00000000;
        rContents[1501] = 8'b00000000;
        rContents[1502] = 8'b00000000;
        rContents[1503] = 8'b00000000;
        rContents[1504] = 8'b00000000;
        rContents[1505] = 8'b00000000;
        rContents[1506] = 8'b00000000;
        rContents[1507] = 8'b00000000;
        rContents[1508] = 8'b00000000;
        rContents[1509] = 8'b00000000;
        rContents[1510] = 8'b00000000;
        rContents[1511] = 8'b00000000;
        rContents[1512] = 8'b00000000;
        rContents[1513] = 8'b00000000;
        rContents[1514] = 8'b00000000;
        rContents[1515] = 8'b00000000;
        rContents[1516] = 8'b00000000;
        rContents[1517] = 8'b00000000;
        rContents[1518] = 8'b00000000;
        rContents[1519] = 8'b00000000;
        rContents[1520] = 8'b00000000;
        rContents[1521] = 8'b00000000;
        rContents[1522] = 8'b00000000;
        rContents[1523] = 8'b00000000;
        rContents[1524] = 8'b00000000;
        rContents[1525] = 8'b00000000;
        rContents[1526] = 8'b00000000;
        rContents[1527] = 8'b00000000;
        rContents[1528] = 8'b00000000;
        rContents[1529] = 8'b00000000;
        rContents[1530] = 8'b00000000;
        rContents[1531] = 8'b00000000;
        rContents[1532] = 8'b00000000;
        rContents[1533] = 8'b00000000;
        rContents[1534] = 8'b00000000;
        rContents[1535] = 8'b00000000;
        rContents[1536] = 8'b01010101;
        rContents[1537] = 8'b10101010;
        rContents[1538] = 8'b01010101;
        rContents[1539] = 8'b11111111;
        rContents[1540] = 8'b11111111;
        rContents[1541] = 8'b00000000;
        rContents[1542] = 8'b11111110;
        rContents[1543] = 8'b10000010;
        rContents[1544] = 8'b00010000;
        rContents[1545] = 8'b10010010;
        rContents[1546] = 8'b11101110;
        rContents[1547] = 8'b00111000;
        rContents[1548] = 8'b00111000;
        rContents[1549] = 8'b01111100;
        rContents[1550] = 8'b00111000;
        rContents[1551] = 8'b10000010;
        rContents[1552] = 8'b10010010;
        rContents[1553] = 8'b11111110;
        rContents[1554] = 8'b10100000;
        rContents[1555] = 8'b10101010;
        rContents[1556] = 8'b00010000;
        rContents[1557] = 8'b01111100;
        rContents[1558] = 8'b00100000;
        rContents[1559] = 8'b00001000;
        rContents[1560] = 8'b11111000;
        rContents[1561] = 8'b00111110;
        rContents[1562] = 8'b01111100;
        rContents[1563] = 8'b00001010;
        rContents[1564] = 8'b00000000;
        rContents[1565] = 8'b01111100;
        rContents[1566] = 8'b00111000;
        rContents[1567] = 8'b00001100;
        rContents[1568] = 8'b00000000;
        rContents[1569] = 8'b00010000;
        rContents[1570] = 8'b00000000;
        rContents[1571] = 8'b11111110;
        rContents[1572] = 8'b00010010;
        rContents[1573] = 8'b01001110;
        rContents[1574] = 8'b01101100;
        rContents[1575] = 8'b00000000;
        rContents[1576] = 8'b00100000;
        rContents[1577] = 8'b00001000;
        rContents[1578] = 8'b00000000;
        rContents[1579] = 8'b00010000;
        rContents[1580] = 8'b00000000;
        rContents[1581] = 8'b00000000;
        rContents[1582] = 8'b00000000;
        rContents[1583] = 8'b01000000;
        rContents[1584] = 8'b10000010;
        rContents[1585] = 8'b00010000;
        rContents[1586] = 8'b01000000;
        rContents[1587] = 8'b00000010;
        rContents[1588] = 8'b00000010;
        rContents[1589] = 8'b00000010;
        rContents[1590] = 8'b10000010;
        rContents[1591] = 8'b00001000;
        rContents[1592] = 8'b10000010;
        rContents[1593] = 8'b00000010;
        rContents[1594] = 8'b00000000;
        rContents[1595] = 8'b00000000;
        rContents[1596] = 8'b00010000;
        rContents[1597] = 8'b11111110;
        rContents[1598] = 8'b00010000;
        rContents[1599] = 8'b00010000;
        rContents[1600] = 8'b10111100;
        rContents[1601] = 8'b01000010;
        rContents[1602] = 8'b10000010;
        rContents[1603] = 8'b10000000;
        rContents[1604] = 8'b10000010;
        rContents[1605] = 8'b10000000;
        rContents[1606] = 8'b10000000;
        rContents[1607] = 8'b10000010;
        rContents[1608] = 8'b10000010;
        rContents[1609] = 8'b00010000;
        rContents[1610] = 8'b00000010;
        rContents[1611] = 8'b10001000;
        rContents[1612] = 8'b10000000;
        rContents[1613] = 8'b10000010;
        rContents[1614] = 8'b10000110;
        rContents[1615] = 8'b10000010;
        rContents[1616] = 8'b10000000;
        rContents[1617] = 8'b10001100;
        rContents[1618] = 8'b10110000;
        rContents[1619] = 8'b00000010;
        rContents[1620] = 8'b00010000;
        rContents[1621] = 8'b10000010;
        rContents[1622] = 8'b00001010;
        rContents[1623] = 8'b10010010;
        rContents[1624] = 8'b01000100;
        rContents[1625] = 8'b00010000;
        rContents[1626] = 8'b01000000;
        rContents[1627] = 8'b00100000;
        rContents[1628] = 8'b00000100;
        rContents[1629] = 8'b00001000;
        rContents[1630] = 8'b00000000;
        rContents[1631] = 8'b00000000;
        rContents[1632] = 8'b00000000;
        rContents[1633] = 8'b11111110;
        rContents[1634] = 8'b10000010;
        rContents[1635] = 8'b10000000;
        rContents[1636] = 8'b10000010;
        rContents[1637] = 8'b11111110;
        rContents[1638] = 8'b10000000;
        rContents[1639] = 8'b10000010;
        rContents[1640] = 8'b10000010;
        rContents[1641] = 8'b00010000;
        rContents[1642] = 8'b00001000;
        rContents[1643] = 8'b11100000;
        rContents[1644] = 8'b00010000;
        rContents[1645] = 8'b10010010;
        rContents[1646] = 8'b10000010;
        rContents[1647] = 8'b10000010;
        rContents[1648] = 8'b10000010;
        rContents[1649] = 8'b10000010;
        rContents[1650] = 8'b10000000;
        rContents[1651] = 8'b11111110;
        rContents[1652] = 8'b10000000;
        rContents[1653] = 8'b10000010;
        rContents[1654] = 8'b00110010;
        rContents[1655] = 8'b10010010;
        rContents[1656] = 8'b00010000;
        rContents[1657] = 8'b10000010;
        rContents[1658] = 8'b00111000;
        rContents[1659] = 8'b00100000;
        rContents[1660] = 8'b00010000;
        rContents[1661] = 8'b00001000;
        rContents[1662] = 8'b00000000;
        rContents[1663] = 8'b00010000;
        rContents[1664] = 8'b00000100;
        rContents[1665] = 8'b11110000;
        rContents[1666] = 8'b00001111;
        rContents[1667] = 8'b11111111;
        rContents[1668] = 8'b11111111;
        rContents[1669] = 8'b00000000;
        rContents[1670] = 8'b00000000;
        rContents[1671] = 8'b11110000;
        rContents[1672] = 8'b00001111;
        rContents[1673] = 8'b11110000;
        rContents[1674] = 8'b00001111;
        rContents[1675] = 8'b00000000;
        rContents[1676] = 8'b11111111;
        rContents[1677] = 8'b00011000;
        rContents[1678] = 8'b11111111;
        rContents[1679] = 8'b11111111;
        rContents[1680] = 8'b11111111;
        rContents[1681] = 8'b11111111;
        rContents[1682] = 8'b11111000;
        rContents[1683] = 8'b11111000;
        rContents[1684] = 8'b00011111;
        rContents[1685] = 8'b00011111;
        rContents[1686] = 8'b11111000;
        rContents[1687] = 8'b00011111;
        rContents[1688] = 8'b00100100;
        rContents[1689] = 8'b00000000;
        rContents[1690] = 8'b00000000;
        rContents[1691] = 8'b00000000;
        rContents[1692] = 8'b00000000;
        rContents[1693] = 8'b00000100;
        rContents[1694] = 8'b00000100;
        rContents[1695] = 8'b00100000;
        rContents[1696] = 8'b00000100;
        rContents[1697] = 8'b00100000;
        rContents[1698] = 8'b01000100;
        rContents[1699] = 8'b01000100;
        rContents[1700] = 8'b10001000;
        rContents[1701] = 8'b11111100;
        rContents[1702] = 8'b01000000;
        rContents[1703] = 8'b00010100;
        rContents[1704] = 8'b00000000;
        rContents[1705] = 8'b00000000;
        rContents[1706] = 8'b00000000;
        rContents[1707] = 8'b00000000;
        rContents[1708] = 8'b00000000;
        rContents[1709] = 8'b00000000;
        rContents[1710] = 8'b00000000;
        rContents[1711] = 8'b00000000;
        rContents[1712] = 8'b00000000;
        rContents[1713] = 8'b00000000;
        rContents[1714] = 8'b00000000;
        rContents[1715] = 8'b00000000;
        rContents[1716] = 8'b00000000;
        rContents[1717] = 8'b00000000;
        rContents[1718] = 8'b00000000;
        rContents[1719] = 8'b00000000;
        rContents[1720] = 8'b00000000;
        rContents[1721] = 8'b00000000;
        rContents[1722] = 8'b00000000;
        rContents[1723] = 8'b00000000;
        rContents[1724] = 8'b00000000;
        rContents[1725] = 8'b00000000;
        rContents[1726] = 8'b00000000;
        rContents[1727] = 8'b00000000;
        rContents[1728] = 8'b00000000;
        rContents[1729] = 8'b00000000;
        rContents[1730] = 8'b00000000;
        rContents[1731] = 8'b00000000;
        rContents[1732] = 8'b00000000;
        rContents[1733] = 8'b00000000;
        rContents[1734] = 8'b00000000;
        rContents[1735] = 8'b00000000;
        rContents[1736] = 8'b00000000;
        rContents[1737] = 8'b00000000;
        rContents[1738] = 8'b00000000;
        rContents[1739] = 8'b00000000;
        rContents[1740] = 8'b00000000;
        rContents[1741] = 8'b00000000;
        rContents[1742] = 8'b00000000;
        rContents[1743] = 8'b00000000;
        rContents[1744] = 8'b00000000;
        rContents[1745] = 8'b00000000;
        rContents[1746] = 8'b00000000;
        rContents[1747] = 8'b00000000;
        rContents[1748] = 8'b00000000;
        rContents[1749] = 8'b00000000;
        rContents[1750] = 8'b00000000;
        rContents[1751] = 8'b00000000;
        rContents[1752] = 8'b00000000;
        rContents[1753] = 8'b00000000;
        rContents[1754] = 8'b00000000;
        rContents[1755] = 8'b00000000;
        rContents[1756] = 8'b00000000;
        rContents[1757] = 8'b00000000;
        rContents[1758] = 8'b00000000;
        rContents[1759] = 8'b00000000;
        rContents[1760] = 8'b00000000;
        rContents[1761] = 8'b00000000;
        rContents[1762] = 8'b00000000;
        rContents[1763] = 8'b00000000;
        rContents[1764] = 8'b00000000;
        rContents[1765] = 8'b00000000;
        rContents[1766] = 8'b00000000;
        rContents[1767] = 8'b00000000;
        rContents[1768] = 8'b00000000;
        rContents[1769] = 8'b00000000;
        rContents[1770] = 8'b00000000;
        rContents[1771] = 8'b00000000;
        rContents[1772] = 8'b00000000;
        rContents[1773] = 8'b00000000;
        rContents[1774] = 8'b00000000;
        rContents[1775] = 8'b00000000;
        rContents[1776] = 8'b00000000;
        rContents[1777] = 8'b00000000;
        rContents[1778] = 8'b00000000;
        rContents[1779] = 8'b00000000;
        rContents[1780] = 8'b00000000;
        rContents[1781] = 8'b00000000;
        rContents[1782] = 8'b00000000;
        rContents[1783] = 8'b00000000;
        rContents[1784] = 8'b00000000;
        rContents[1785] = 8'b00000000;
        rContents[1786] = 8'b00000000;
        rContents[1787] = 8'b00000000;
        rContents[1788] = 8'b00000000;
        rContents[1789] = 8'b00000000;
        rContents[1790] = 8'b00000000;
        rContents[1791] = 8'b00000000;
        rContents[1792] = 8'b01010101;
        rContents[1793] = 8'b10101010;
        rContents[1794] = 8'b11111111;
        rContents[1795] = 8'b10101010;
        rContents[1796] = 8'b11111111;
        rContents[1797] = 8'b00000000;
        rContents[1798] = 8'b11111110;
        rContents[1799] = 8'b10000010;
        rContents[1800] = 8'b00010000;
        rContents[1801] = 8'b10000010;
        rContents[1802] = 8'b11111110;
        rContents[1803] = 8'b00111000;
        rContents[1804] = 8'b00111000;
        rContents[1805] = 8'b00111000;
        rContents[1806] = 8'b00010000;
        rContents[1807] = 8'b10000010;
        rContents[1808] = 8'b10000010;
        rContents[1809] = 8'b11111110;
        rContents[1810] = 8'b10100000;
        rContents[1811] = 8'b10101010;
        rContents[1812] = 8'b00010000;
        rContents[1813] = 8'b00111000;
        rContents[1814] = 8'b00000000;
        rContents[1815] = 8'b00000000;
        rContents[1816] = 8'b11110000;
        rContents[1817] = 8'b00011110;
        rContents[1818] = 8'b00111000;
        rContents[1819] = 8'b00001010;
        rContents[1820] = 8'b00000000;
        rContents[1821] = 8'b00111000;
        rContents[1822] = 8'b00010000;
        rContents[1823] = 8'b00000100;
        rContents[1824] = 8'b00000000;
        rContents[1825] = 8'b00000000;
        rContents[1826] = 8'b00000000;
        rContents[1827] = 8'b01000100;
        rContents[1828] = 8'b11111110;
        rContents[1829] = 8'b10001010;
        rContents[1830] = 8'b10000010;
        rContents[1831] = 8'b00000000;
        rContents[1832] = 8'b00010000;
        rContents[1833] = 8'b00010000;
        rContents[1834] = 8'b00000000;
        rContents[1835] = 8'b00010000;
        rContents[1836] = 8'b00000000;
        rContents[1837] = 8'b00000000;
        rContents[1838] = 8'b00000000;
        rContents[1839] = 8'b10000000;
        rContents[1840] = 8'b10000010;
        rContents[1841] = 8'b00010000;
        rContents[1842] = 8'b10000000;
        rContents[1843] = 8'b10000010;
        rContents[1844] = 8'b00000010;
        rContents[1845] = 8'b00000010;
        rContents[1846] = 8'b10000010;
        rContents[1847] = 8'b00010000;
        rContents[1848] = 8'b10000010;
        rContents[1849] = 8'b00000010;
        rContents[1850] = 8'b00010000;
        rContents[1851] = 8'b00010000;
        rContents[1852] = 8'b00001100;
        rContents[1853] = 8'b00000000;
        rContents[1854] = 8'b01100000;
        rContents[1855] = 8'b00000000;
        rContents[1856] = 8'b10000000;
        rContents[1857] = 8'b01000010;
        rContents[1858] = 8'b10000010;
        rContents[1859] = 8'b10000000;
        rContents[1860] = 8'b10000010;
        rContents[1861] = 8'b10000000;
        rContents[1862] = 8'b10000000;
        rContents[1863] = 8'b10000010;
        rContents[1864] = 8'b10000010;
        rContents[1865] = 8'b00010000;
        rContents[1866] = 8'b00000010;
        rContents[1867] = 8'b10000100;
        rContents[1868] = 8'b10000000;
        rContents[1869] = 8'b10000010;
        rContents[1870] = 8'b10000010;
        rContents[1871] = 8'b10000010;
        rContents[1872] = 8'b10000000;
        rContents[1873] = 8'b10001100;
        rContents[1874] = 8'b10001100;
        rContents[1875] = 8'b00000010;
        rContents[1876] = 8'b00010000;
        rContents[1877] = 8'b10000010;
        rContents[1878] = 8'b00001010;
        rContents[1879] = 8'b10010010;
        rContents[1880] = 8'b10000010;
        rContents[1881] = 8'b00010000;
        rContents[1882] = 8'b10000000;
        rContents[1883] = 8'b00100000;
        rContents[1884] = 8'b00000010;
        rContents[1885] = 8'b00001000;
        rContents[1886] = 8'b00000000;
        rContents[1887] = 8'b00000000;
        rContents[1888] = 8'b00000000;
        rContents[1889] = 8'b10000010;
        rContents[1890] = 8'b10000010;
        rContents[1891] = 8'b10000000;
        rContents[1892] = 8'b10000010;
        rContents[1893] = 8'b10000000;
        rContents[1894] = 8'b10000000;
        rContents[1895] = 8'b10000010;
        rContents[1896] = 8'b10000010;
        rContents[1897] = 8'b00010000;
        rContents[1898] = 8'b00001000;
        rContents[1899] = 8'b10011000;
        rContents[1900] = 8'b00010000;
        rContents[1901] = 8'b10000010;
        rContents[1902] = 8'b10000010;
        rContents[1903] = 8'b10000010;
        rContents[1904] = 8'b10000010;
        rContents[1905] = 8'b10000010;
        rContents[1906] = 8'b10000000;
        rContents[1907] = 8'b00000010;
        rContents[1908] = 8'b10000000;
        rContents[1909] = 8'b10000010;
        rContents[1910] = 8'b00001010;
        rContents[1911] = 8'b10010010;
        rContents[1912] = 8'b00101000;
        rContents[1913] = 8'b10000010;
        rContents[1914] = 8'b01000000;
        rContents[1915] = 8'b00100000;
        rContents[1916] = 8'b00010000;
        rContents[1917] = 8'b00001000;
        rContents[1918] = 8'b00000000;
        rContents[1919] = 8'b00010000;
        rContents[1920] = 8'b00000100;
        rContents[1921] = 8'b11110000;
        rContents[1922] = 8'b00001111;
        rContents[1923] = 8'b11111111;
        rContents[1924] = 8'b11111111;
        rContents[1925] = 8'b00000000;
        rContents[1926] = 8'b00000000;
        rContents[1927] = 8'b11110000;
        rContents[1928] = 8'b00001111;
        rContents[1929] = 8'b11110000;
        rContents[1930] = 8'b00001111;
        rContents[1931] = 8'b00000000;
        rContents[1932] = 8'b11111111;
        rContents[1933] = 8'b00011000;
        rContents[1934] = 8'b00000000;
        rContents[1935] = 8'b00011000;
        rContents[1936] = 8'b00000000;
        rContents[1937] = 8'b00011000;
        rContents[1938] = 8'b00011000;
        rContents[1939] = 8'b00000000;
        rContents[1940] = 8'b00011000;
        rContents[1941] = 8'b00000000;
        rContents[1942] = 8'b00011000;
        rContents[1943] = 8'b00011000;
        rContents[1944] = 8'b00100100;
        rContents[1945] = 8'b11111111;
        rContents[1946] = 8'b11100111;
        rContents[1947] = 8'b11111111;
        rContents[1948] = 8'b11100111;
        rContents[1949] = 8'b11100100;
        rContents[1950] = 8'b11111100;
        rContents[1951] = 8'b00100111;
        rContents[1952] = 8'b11100100;
        rContents[1953] = 8'b00100111;
        rContents[1954] = 8'b00101000;
        rContents[1955] = 8'b01000100;
        rContents[1956] = 8'b10001100;
        rContents[1957] = 8'b10000000;
        rContents[1958] = 8'b10000010;
        rContents[1959] = 8'b00010100;
        rContents[1960] = 8'b00000000;
        rContents[1961] = 8'b00000000;
        rContents[1962] = 8'b00000000;
        rContents[1963] = 8'b00000000;
        rContents[1964] = 8'b00000000;
        rContents[1965] = 8'b00000000;
        rContents[1966] = 8'b00000000;
        rContents[1967] = 8'b00000000;
        rContents[1968] = 8'b00000000;
        rContents[1969] = 8'b00000000;
        rContents[1970] = 8'b00000000;
        rContents[1971] = 8'b00000000;
        rContents[1972] = 8'b00000000;
        rContents[1973] = 8'b00000000;
        rContents[1974] = 8'b00000000;
        rContents[1975] = 8'b00000000;
        rContents[1976] = 8'b00000000;
        rContents[1977] = 8'b00000000;
        rContents[1978] = 8'b00000000;
        rContents[1979] = 8'b00000000;
        rContents[1980] = 8'b00000000;
        rContents[1981] = 8'b00000000;
        rContents[1982] = 8'b00000000;
        rContents[1983] = 8'b00000000;
        rContents[1984] = 8'b00000000;
        rContents[1985] = 8'b00000000;
        rContents[1986] = 8'b00000000;
        rContents[1987] = 8'b00000000;
        rContents[1988] = 8'b00000000;
        rContents[1989] = 8'b00000000;
        rContents[1990] = 8'b00000000;
        rContents[1991] = 8'b00000000;
        rContents[1992] = 8'b00000000;
        rContents[1993] = 8'b00000000;
        rContents[1994] = 8'b00000000;
        rContents[1995] = 8'b00000000;
        rContents[1996] = 8'b00000000;
        rContents[1997] = 8'b00000000;
        rContents[1998] = 8'b00000000;
        rContents[1999] = 8'b00000000;
        rContents[2000] = 8'b00000000;
        rContents[2001] = 8'b00000000;
        rContents[2002] = 8'b00000000;
        rContents[2003] = 8'b00000000;
        rContents[2004] = 8'b00000000;
        rContents[2005] = 8'b00000000;
        rContents[2006] = 8'b00000000;
        rContents[2007] = 8'b00000000;
        rContents[2008] = 8'b00000000;
        rContents[2009] = 8'b00000000;
        rContents[2010] = 8'b00000000;
        rContents[2011] = 8'b00000000;
        rContents[2012] = 8'b00000000;
        rContents[2013] = 8'b00000000;
        rContents[2014] = 8'b00000000;
        rContents[2015] = 8'b00000000;
        rContents[2016] = 8'b00000000;
        rContents[2017] = 8'b00000000;
        rContents[2018] = 8'b00000000;
        rContents[2019] = 8'b00000000;
        rContents[2020] = 8'b00000000;
        rContents[2021] = 8'b00000000;
        rContents[2022] = 8'b00000000;
        rContents[2023] = 8'b00000000;
        rContents[2024] = 8'b00000000;
        rContents[2025] = 8'b00000000;
        rContents[2026] = 8'b00000000;
        rContents[2027] = 8'b00000000;
        rContents[2028] = 8'b00000000;
        rContents[2029] = 8'b00000000;
        rContents[2030] = 8'b00000000;
        rContents[2031] = 8'b00000000;
        rContents[2032] = 8'b00000000;
        rContents[2033] = 8'b00000000;
        rContents[2034] = 8'b00000000;
        rContents[2035] = 8'b00000000;
        rContents[2036] = 8'b00000000;
        rContents[2037] = 8'b00000000;
        rContents[2038] = 8'b00000000;
        rContents[2039] = 8'b00000000;
        rContents[2040] = 8'b00000000;
        rContents[2041] = 8'b00000000;
        rContents[2042] = 8'b00000000;
        rContents[2043] = 8'b00000000;
        rContents[2044] = 8'b00000000;
        rContents[2045] = 8'b00000000;
        rContents[2046] = 8'b00000000;
        rContents[2047] = 8'b00000000;
        rContents[2048] = 8'b01010101;
        rContents[2049] = 8'b10101010;
        rContents[2050] = 8'b01010101;
        rContents[2051] = 8'b11111111;
        rContents[2052] = 8'b11111111;
        rContents[2053] = 8'b00000000;
        rContents[2054] = 8'b11111110;
        rContents[2055] = 8'b11111110;
        rContents[2056] = 8'b00111000;
        rContents[2057] = 8'b01111100;
        rContents[2058] = 8'b01111100;
        rContents[2059] = 8'b00010000;
        rContents[2060] = 8'b00010000;
        rContents[2061] = 8'b11111110;
        rContents[2062] = 8'b11111110;
        rContents[2063] = 8'b11111110;
        rContents[2064] = 8'b11111110;
        rContents[2065] = 8'b11111110;
        rContents[2066] = 8'b01100000;
        rContents[2067] = 8'b01100110;
        rContents[2068] = 8'b00010000;
        rContents[2069] = 8'b00010000;
        rContents[2070] = 8'b00000000;
        rContents[2071] = 8'b00000000;
        rContents[2072] = 8'b11000000;
        rContents[2073] = 8'b00000110;
        rContents[2074] = 8'b00010000;
        rContents[2075] = 8'b00001010;
        rContents[2076] = 8'b00000000;
        rContents[2077] = 8'b00010000;
        rContents[2078] = 8'b11111110;
        rContents[2079] = 8'b01111100;
        rContents[2080] = 8'b00000000;
        rContents[2081] = 8'b00010000;
        rContents[2082] = 8'b00000000;
        rContents[2083] = 8'b01000100;
        rContents[2084] = 8'b00010000;
        rContents[2085] = 8'b10001110;
        rContents[2086] = 8'b10000010;
        rContents[2087] = 8'b00000000;
        rContents[2088] = 8'b00001000;
        rContents[2089] = 8'b00100000;
        rContents[2090] = 8'b00000000;
        rContents[2091] = 8'b00010000;
        rContents[2092] = 8'b00010000;
        rContents[2093] = 8'b00000000;
        rContents[2094] = 8'b00010000;
        rContents[2095] = 8'b10000000;
        rContents[2096] = 8'b01111100;
        rContents[2097] = 8'b00111000;
        rContents[2098] = 8'b11111110;
        rContents[2099] = 8'b01111100;
        rContents[2100] = 8'b00000010;
        rContents[2101] = 8'b11111100;
        rContents[2102] = 8'b01111100;
        rContents[2103] = 8'b00010000;
        rContents[2104] = 8'b01111100;
        rContents[2105] = 8'b00000010;
        rContents[2106] = 8'b00000000;
        rContents[2107] = 8'b00010000;
        rContents[2108] = 8'b00000010;
        rContents[2109] = 8'b00000000;
        rContents[2110] = 8'b10000000;
        rContents[2111] = 8'b00010000;
        rContents[2112] = 8'b11111110;
        rContents[2113] = 8'b10000010;
        rContents[2114] = 8'b11111110;
        rContents[2115] = 8'b11111110;
        rContents[2116] = 8'b11111110;
        rContents[2117] = 8'b11111110;
        rContents[2118] = 8'b10000000;
        rContents[2119] = 8'b11111110;
        rContents[2120] = 8'b10000010;
        rContents[2121] = 8'b11111110;
        rContents[2122] = 8'b11111110;
        rContents[2123] = 8'b10000010;
        rContents[2124] = 8'b11111110;
        rContents[2125] = 8'b10000010;
        rContents[2126] = 8'b10000010;
        rContents[2127] = 8'b11111110;
        rContents[2128] = 8'b10000000;
        rContents[2129] = 8'b11110010;
        rContents[2130] = 8'b10000010;
        rContents[2131] = 8'b11111110;
        rContents[2132] = 8'b00010000;
        rContents[2133] = 8'b11111110;
        rContents[2134] = 8'b00000110;
        rContents[2135] = 8'b11111110;
        rContents[2136] = 8'b10000010;
        rContents[2137] = 8'b00010000;
        rContents[2138] = 8'b11111110;
        rContents[2139] = 8'b00111000;
        rContents[2140] = 8'b00000010;
        rContents[2141] = 8'b00111000;
        rContents[2142] = 8'b00000000;
        rContents[2143] = 8'b11111110;
        rContents[2144] = 8'b00000000;
        rContents[2145] = 8'b11111110;
        rContents[2146] = 8'b11111110;
        rContents[2147] = 8'b11111110;
        rContents[2148] = 8'b11111110;
        rContents[2149] = 8'b11111110;
        rContents[2150] = 8'b10000000;
        rContents[2151] = 8'b11111110;
        rContents[2152] = 8'b10000010;
        rContents[2153] = 8'b00010000;
        rContents[2154] = 8'b00001000;
        rContents[2155] = 8'b10000110;
        rContents[2156] = 8'b00010000;
        rContents[2157] = 8'b10000010;
        rContents[2158] = 8'b10000010;
        rContents[2159] = 8'b11111110;
        rContents[2160] = 8'b11111110;
        rContents[2161] = 8'b11111110;
        rContents[2162] = 8'b10000000;
        rContents[2163] = 8'b11111110;
        rContents[2164] = 8'b11111110;
        rContents[2165] = 8'b11111110;
        rContents[2166] = 8'b00000110;
        rContents[2167] = 8'b11111110;
        rContents[2168] = 8'b11000110;
        rContents[2169] = 8'b11111110;
        rContents[2170] = 8'b11111110;
        rContents[2171] = 8'b00011000;
        rContents[2172] = 8'b00010000;
        rContents[2173] = 8'b00110000;
        rContents[2174] = 8'b00000000;
        rContents[2175] = 8'b00010000;
        rContents[2176] = 8'b01111100;
        rContents[2177] = 8'b11110000;
        rContents[2178] = 8'b00001111;
        rContents[2179] = 8'b11111111;
        rContents[2180] = 8'b11111111;
        rContents[2181] = 8'b00000000;
        rContents[2182] = 8'b00000000;
        rContents[2183] = 8'b11110000;
        rContents[2184] = 8'b00001111;
        rContents[2185] = 8'b11110000;
        rContents[2186] = 8'b00001111;
        rContents[2187] = 8'b00000000;
        rContents[2188] = 8'b11111111;
        rContents[2189] = 8'b00011000;
        rContents[2190] = 8'b00000000;
        rContents[2191] = 8'b00011000;
        rContents[2192] = 8'b00000000;
        rContents[2193] = 8'b00011000;
        rContents[2194] = 8'b00011000;
        rContents[2195] = 8'b00000000;
        rContents[2196] = 8'b00011000;
        rContents[2197] = 8'b00000000;
        rContents[2198] = 8'b00011000;
        rContents[2199] = 8'b00011000;
        rContents[2200] = 8'b00100100;
        rContents[2201] = 8'b00000000;
        rContents[2202] = 8'b00100100;
        rContents[2203] = 8'b00000000;
        rContents[2204] = 8'b00100100;
        rContents[2205] = 8'b00100100;
        rContents[2206] = 8'b00000000;
        rContents[2207] = 8'b00100100;
        rContents[2208] = 8'b00100100;
        rContents[2209] = 8'b00100100;
        rContents[2210] = 8'b11101110;
        rContents[2211] = 8'b01000100;
        rContents[2212] = 8'b01110010;
        rContents[2213] = 8'b10000000;
        rContents[2214] = 8'b11111110;
        rContents[2215] = 8'b00001100;
        rContents[2216] = 8'b00000000;
        rContents[2217] = 8'b00000000;
        rContents[2218] = 8'b00000000;
        rContents[2219] = 8'b00000000;
        rContents[2220] = 8'b00000000;
        rContents[2221] = 8'b00000000;
        rContents[2222] = 8'b00000000;
        rContents[2223] = 8'b00000000;
        rContents[2224] = 8'b00000000;
        rContents[2225] = 8'b00000000;
        rContents[2226] = 8'b00000000;
        rContents[2227] = 8'b00000000;
        rContents[2228] = 8'b00000000;
        rContents[2229] = 8'b00000000;
        rContents[2230] = 8'b00000000;
        rContents[2231] = 8'b00000000;
        rContents[2232] = 8'b00000000;
        rContents[2233] = 8'b00000000;
        rContents[2234] = 8'b00000000;
        rContents[2235] = 8'b00000000;
        rContents[2236] = 8'b00000000;
        rContents[2237] = 8'b00000000;
        rContents[2238] = 8'b00000000;
        rContents[2239] = 8'b00000000;
        rContents[2240] = 8'b00000000;
        rContents[2241] = 8'b00000000;
        rContents[2242] = 8'b00000000;
        rContents[2243] = 8'b00000000;
        rContents[2244] = 8'b00000000;
        rContents[2245] = 8'b00000000;
        rContents[2246] = 8'b00000000;
        rContents[2247] = 8'b00000000;
        rContents[2248] = 8'b00000000;
        rContents[2249] = 8'b00000000;
        rContents[2250] = 8'b00000000;
        rContents[2251] = 8'b00000000;
        rContents[2252] = 8'b00000000;
        rContents[2253] = 8'b00000000;
        rContents[2254] = 8'b00000000;
        rContents[2255] = 8'b00000000;
        rContents[2256] = 8'b00000000;
        rContents[2257] = 8'b00000000;
        rContents[2258] = 8'b00000000;
        rContents[2259] = 8'b00000000;
        rContents[2260] = 8'b00000000;
        rContents[2261] = 8'b00000000;
        rContents[2262] = 8'b00000000;
        rContents[2263] = 8'b00000000;
        rContents[2264] = 8'b00000000;
        rContents[2265] = 8'b00000000;
        rContents[2266] = 8'b00000000;
        rContents[2267] = 8'b00000000;
        rContents[2268] = 8'b00000000;
        rContents[2269] = 8'b00000000;
        rContents[2270] = 8'b00000000;
        rContents[2271] = 8'b00000000;
        rContents[2272] = 8'b00000000;
        rContents[2273] = 8'b00000000;
        rContents[2274] = 8'b00000000;
        rContents[2275] = 8'b00000000;
        rContents[2276] = 8'b00000000;
        rContents[2277] = 8'b00000000;
        rContents[2278] = 8'b00000000;
        rContents[2279] = 8'b00000000;
        rContents[2280] = 8'b00000000;
        rContents[2281] = 8'b00000000;
        rContents[2282] = 8'b00000000;
        rContents[2283] = 8'b00000000;
        rContents[2284] = 8'b00000000;
        rContents[2285] = 8'b00000000;
        rContents[2286] = 8'b00000000;
        rContents[2287] = 8'b00000000;
        rContents[2288] = 8'b00000000;
        rContents[2289] = 8'b00000000;
        rContents[2290] = 8'b00000000;
        rContents[2291] = 8'b00000000;
        rContents[2292] = 8'b00000000;
        rContents[2293] = 8'b00000000;
        rContents[2294] = 8'b00000000;
        rContents[2295] = 8'b00000000;
        rContents[2296] = 8'b00000000;
        rContents[2297] = 8'b00000000;
        rContents[2298] = 8'b00000000;
        rContents[2299] = 8'b00000000;
        rContents[2300] = 8'b00000000;
        rContents[2301] = 8'b00000000;
        rContents[2302] = 8'b00000000;
        rContents[2303] = 8'b00000000;
        rContents[2304] = 8'b01010101;
        rContents[2305] = 8'b10101010;
        rContents[2306] = 8'b11111111;
        rContents[2307] = 8'b10101010;
        rContents[2308] = 8'b11111111;
        rContents[2309] = 8'b00000000;
        rContents[2310] = 8'b00000000;
        rContents[2311] = 8'b00000000;
        rContents[2312] = 8'b00000000;
        rContents[2313] = 8'b00000000;
        rContents[2314] = 8'b00000000;
        rContents[2315] = 8'b00000000;
        rContents[2316] = 8'b00000000;
        rContents[2317] = 8'b00000000;
        rContents[2318] = 8'b00000000;
        rContents[2319] = 8'b00000000;
        rContents[2320] = 8'b00000000;
        rContents[2321] = 8'b00000000;
        rContents[2322] = 8'b00000000;
        rContents[2323] = 8'b00000000;
        rContents[2324] = 8'b00000000;
        rContents[2325] = 8'b00000000;
        rContents[2326] = 8'b00000000;
        rContents[2327] = 8'b00000000;
        rContents[2328] = 8'b00000000;
        rContents[2329] = 8'b00000000;
        rContents[2330] = 8'b00000000;
        rContents[2331] = 8'b00000000;
        rContents[2332] = 8'b00000000;
        rContents[2333] = 8'b00000000;
        rContents[2334] = 8'b00000000;
        rContents[2335] = 8'b00000000;
        rContents[2336] = 8'b00000000;
        rContents[2337] = 8'b00000000;
        rContents[2338] = 8'b00000000;
        rContents[2339] = 8'b00000000;
        rContents[2340] = 8'b00000000;
        rContents[2341] = 8'b00000000;
        rContents[2342] = 8'b00000000;
        rContents[2343] = 8'b00000000;
        rContents[2344] = 8'b00000000;
        rContents[2345] = 8'b00000000;
        rContents[2346] = 8'b00000000;
        rContents[2347] = 8'b00000000;
        rContents[2348] = 8'b00100000;
        rContents[2349] = 8'b00000000;
        rContents[2350] = 8'b00000000;
        rContents[2351] = 8'b00000000;
        rContents[2352] = 8'b00000000;
        rContents[2353] = 8'b00000000;
        rContents[2354] = 8'b00000000;
        rContents[2355] = 8'b00000000;
        rContents[2356] = 8'b00000000;
        rContents[2357] = 8'b00000000;
        rContents[2358] = 8'b00000000;
        rContents[2359] = 8'b00000000;
        rContents[2360] = 8'b00000000;
        rContents[2361] = 8'b00000000;
        rContents[2362] = 8'b00000000;
        rContents[2363] = 8'b00100000;
        rContents[2364] = 8'b00000000;
        rContents[2365] = 8'b00000000;
        rContents[2366] = 8'b00000000;
        rContents[2367] = 8'b00000000;
        rContents[2368] = 8'b00000000;
        rContents[2369] = 8'b00000000;
        rContents[2370] = 8'b00000000;
        rContents[2371] = 8'b00000000;
        rContents[2372] = 8'b00000000;
        rContents[2373] = 8'b00000000;
        rContents[2374] = 8'b00000000;
        rContents[2375] = 8'b00000000;
        rContents[2376] = 8'b00000000;
        rContents[2377] = 8'b00000000;
        rContents[2378] = 8'b00000000;
        rContents[2379] = 8'b00000000;
        rContents[2380] = 8'b00000000;
        rContents[2381] = 8'b00000000;
        rContents[2382] = 8'b00000000;
        rContents[2383] = 8'b00000000;
        rContents[2384] = 8'b00000000;
        rContents[2385] = 8'b00000000;
        rContents[2386] = 8'b00000000;
        rContents[2387] = 8'b00000000;
        rContents[2388] = 8'b00000000;
        rContents[2389] = 8'b00000000;
        rContents[2390] = 8'b00000000;
        rContents[2391] = 8'b00000000;
        rContents[2392] = 8'b00000000;
        rContents[2393] = 8'b00000000;
        rContents[2394] = 8'b00000000;
        rContents[2395] = 8'b00000000;
        rContents[2396] = 8'b00000000;
        rContents[2397] = 8'b00000000;
        rContents[2398] = 8'b00000000;
        rContents[2399] = 8'b00000000;
        rContents[2400] = 8'b00000000;
        rContents[2401] = 8'b00000000;
        rContents[2402] = 8'b00000000;
        rContents[2403] = 8'b00000000;
        rContents[2404] = 8'b00000000;
        rContents[2405] = 8'b00000000;
        rContents[2406] = 8'b00000000;
        rContents[2407] = 8'b00000010;
        rContents[2408] = 8'b00000000;
        rContents[2409] = 8'b00000000;
        rContents[2410] = 8'b00110000;
        rContents[2411] = 8'b00000000;
        rContents[2412] = 8'b00000000;
        rContents[2413] = 8'b00000000;
        rContents[2414] = 8'b00000000;
        rContents[2415] = 8'b00000000;
        rContents[2416] = 8'b10000000;
        rContents[2417] = 8'b00000010;
        rContents[2418] = 8'b00000000;
        rContents[2419] = 8'b00000000;
        rContents[2420] = 8'b00000000;
        rContents[2421] = 8'b00000000;
        rContents[2422] = 8'b00000000;
        rContents[2423] = 8'b00000000;
        rContents[2424] = 8'b00000000;
        rContents[2425] = 8'b00000010;
        rContents[2426] = 8'b00000000;
        rContents[2427] = 8'b00000000;
        rContents[2428] = 8'b00000000;
        rContents[2429] = 8'b00000000;
        rContents[2430] = 8'b00000000;
        rContents[2431] = 8'b00000000;
        rContents[2432] = 8'b00000000;
        rContents[2433] = 8'b11110000;
        rContents[2434] = 8'b00001111;
        rContents[2435] = 8'b11111111;
        rContents[2436] = 8'b11111111;
        rContents[2437] = 8'b00000000;
        rContents[2438] = 8'b00000000;
        rContents[2439] = 8'b11110000;
        rContents[2440] = 8'b00001111;
        rContents[2441] = 8'b11110000;
        rContents[2442] = 8'b00001111;
        rContents[2443] = 8'b00000000;
        rContents[2444] = 8'b11111111;
        rContents[2445] = 8'b00011000;
        rContents[2446] = 8'b00000000;
        rContents[2447] = 8'b00011000;
        rContents[2448] = 8'b00000000;
        rContents[2449] = 8'b00011000;
        rContents[2450] = 8'b00011000;
        rContents[2451] = 8'b00000000;
        rContents[2452] = 8'b00011000;
        rContents[2453] = 8'b00000000;
        rContents[2454] = 8'b00011000;
        rContents[2455] = 8'b00011000;
        rContents[2456] = 8'b00100100;
        rContents[2457] = 8'b00000000;
        rContents[2458] = 8'b00100100;
        rContents[2459] = 8'b00000000;
        rContents[2460] = 8'b00100100;
        rContents[2461] = 8'b00100100;
        rContents[2462] = 8'b00000000;
        rContents[2463] = 8'b00100100;
        rContents[2464] = 8'b00100100;
        rContents[2465] = 8'b00100100;
        rContents[2466] = 8'b00000000;
        rContents[2467] = 8'b00000000;
        rContents[2468] = 8'b00000000;
        rContents[2469] = 8'b00000000;
        rContents[2470] = 8'b00000000;
        rContents[2471] = 8'b00000000;
        rContents[2472] = 8'b00000000;
        rContents[2473] = 8'b00000000;
        rContents[2474] = 8'b00000000;
        rContents[2475] = 8'b00000000;
        rContents[2476] = 8'b00000000;
        rContents[2477] = 8'b00000000;
        rContents[2478] = 8'b00000000;
        rContents[2479] = 8'b00000000;
        rContents[2480] = 8'b00000000;
        rContents[2481] = 8'b00000000;
        rContents[2482] = 8'b00000000;
        rContents[2483] = 8'b00000000;
        rContents[2484] = 8'b00000000;
        rContents[2485] = 8'b00000000;
        rContents[2486] = 8'b00000000;
        rContents[2487] = 8'b00000000;
        rContents[2488] = 8'b00000000;
        rContents[2489] = 8'b00000000;
        rContents[2490] = 8'b00000000;
        rContents[2491] = 8'b00000000;
        rContents[2492] = 8'b00000000;
        rContents[2493] = 8'b00000000;
        rContents[2494] = 8'b00000000;
        rContents[2495] = 8'b00000000;
        rContents[2496] = 8'b00000000;
        rContents[2497] = 8'b00000000;
        rContents[2498] = 8'b00000000;
        rContents[2499] = 8'b00000000;
        rContents[2500] = 8'b00000000;
        rContents[2501] = 8'b00000000;
        rContents[2502] = 8'b00000000;
        rContents[2503] = 8'b00000000;
        rContents[2504] = 8'b00000000;
        rContents[2505] = 8'b00000000;
        rContents[2506] = 8'b00000000;
        rContents[2507] = 8'b00000000;
        rContents[2508] = 8'b00000000;
        rContents[2509] = 8'b00000000;
        rContents[2510] = 8'b00000000;
        rContents[2511] = 8'b00000000;
        rContents[2512] = 8'b00000000;
        rContents[2513] = 8'b00000000;
        rContents[2514] = 8'b00000000;
        rContents[2515] = 8'b00000000;
        rContents[2516] = 8'b00000000;
        rContents[2517] = 8'b00000000;
        rContents[2518] = 8'b00000000;
        rContents[2519] = 8'b00000000;
        rContents[2520] = 8'b00000000;
        rContents[2521] = 8'b00000000;
        rContents[2522] = 8'b00000000;
        rContents[2523] = 8'b00000000;
        rContents[2524] = 8'b00000000;
        rContents[2525] = 8'b00000000;
        rContents[2526] = 8'b00000000;
        rContents[2527] = 8'b00000000;
        rContents[2528] = 8'b00000000;
        rContents[2529] = 8'b00000000;
        rContents[2530] = 8'b00000000;
        rContents[2531] = 8'b00000000;
        rContents[2532] = 8'b00000000;
        rContents[2533] = 8'b00000000;
        rContents[2534] = 8'b00000000;
        rContents[2535] = 8'b00000000;
        rContents[2536] = 8'b00000000;
        rContents[2537] = 8'b00000000;
        rContents[2538] = 8'b00000000;
        rContents[2539] = 8'b00000000;
        rContents[2540] = 8'b00000000;
        rContents[2541] = 8'b00000000;
        rContents[2542] = 8'b00000000;
        rContents[2543] = 8'b00000000;
        rContents[2544] = 8'b00000000;
        rContents[2545] = 8'b00000000;
        rContents[2546] = 8'b00000000;
        rContents[2547] = 8'b00000000;
        rContents[2548] = 8'b00000000;
        rContents[2549] = 8'b00000000;
        rContents[2550] = 8'b00000000;
        rContents[2551] = 8'b00000000;
        rContents[2552] = 8'b00000000;
        rContents[2553] = 8'b00000000;
        rContents[2554] = 8'b00000000;
        rContents[2555] = 8'b00000000;
        rContents[2556] = 8'b00000000;
        rContents[2557] = 8'b00000000;
        rContents[2558] = 8'b00000000;
        rContents[2559] = 8'b00000000;
        rContents[2560] = 8'b01010101;
        rContents[2561] = 8'b10101010;
        rContents[2562] = 8'b01010101;
        rContents[2563] = 8'b11111111;
        rContents[2564] = 8'b11111111;
        rContents[2565] = 8'b00000000;
        rContents[2566] = 8'b00000000;
        rContents[2567] = 8'b00000000;
        rContents[2568] = 8'b00000000;
        rContents[2569] = 8'b00000000;
        rContents[2570] = 8'b00000000;
        rContents[2571] = 8'b00000000;
        rContents[2572] = 8'b00000000;
        rContents[2573] = 8'b00000000;
        rContents[2574] = 8'b00000000;
        rContents[2575] = 8'b00000000;
        rContents[2576] = 8'b00000000;
        rContents[2577] = 8'b00000000;
        rContents[2578] = 8'b00000000;
        rContents[2579] = 8'b00000000;
        rContents[2580] = 8'b00000000;
        rContents[2581] = 8'b00000000;
        rContents[2582] = 8'b00000000;
        rContents[2583] = 8'b00000000;
        rContents[2584] = 8'b00000000;
        rContents[2585] = 8'b00000000;
        rContents[2586] = 8'b00000000;
        rContents[2587] = 8'b00000000;
        rContents[2588] = 8'b00000000;
        rContents[2589] = 8'b00000000;
        rContents[2590] = 8'b00000000;
        rContents[2591] = 8'b00000000;
        rContents[2592] = 8'b00000000;
        rContents[2593] = 8'b00000000;
        rContents[2594] = 8'b00000000;
        rContents[2595] = 8'b00000000;
        rContents[2596] = 8'b00000000;
        rContents[2597] = 8'b00000000;
        rContents[2598] = 8'b00000000;
        rContents[2599] = 8'b00000000;
        rContents[2600] = 8'b00000000;
        rContents[2601] = 8'b00000000;
        rContents[2602] = 8'b00000000;
        rContents[2603] = 8'b00000000;
        rContents[2604] = 8'b00000000;
        rContents[2605] = 8'b00000000;
        rContents[2606] = 8'b00000000;
        rContents[2607] = 8'b00000000;
        rContents[2608] = 8'b00000000;
        rContents[2609] = 8'b00000000;
        rContents[2610] = 8'b00000000;
        rContents[2611] = 8'b00000000;
        rContents[2612] = 8'b00000000;
        rContents[2613] = 8'b00000000;
        rContents[2614] = 8'b00000000;
        rContents[2615] = 8'b00000000;
        rContents[2616] = 8'b00000000;
        rContents[2617] = 8'b00000000;
        rContents[2618] = 8'b00000000;
        rContents[2619] = 8'b00000000;
        rContents[2620] = 8'b00000000;
        rContents[2621] = 8'b00000000;
        rContents[2622] = 8'b00000000;
        rContents[2623] = 8'b00000000;
        rContents[2624] = 8'b00000000;
        rContents[2625] = 8'b00000000;
        rContents[2626] = 8'b00000000;
        rContents[2627] = 8'b00000000;
        rContents[2628] = 8'b00000000;
        rContents[2629] = 8'b00000000;
        rContents[2630] = 8'b00000000;
        rContents[2631] = 8'b00000000;
        rContents[2632] = 8'b00000000;
        rContents[2633] = 8'b00000000;
        rContents[2634] = 8'b00000000;
        rContents[2635] = 8'b00000000;
        rContents[2636] = 8'b00000000;
        rContents[2637] = 8'b00000000;
        rContents[2638] = 8'b00000000;
        rContents[2639] = 8'b00000000;
        rContents[2640] = 8'b00000000;
        rContents[2641] = 8'b00000000;
        rContents[2642] = 8'b00000000;
        rContents[2643] = 8'b00000000;
        rContents[2644] = 8'b00000000;
        rContents[2645] = 8'b00000000;
        rContents[2646] = 8'b00000000;
        rContents[2647] = 8'b00000000;
        rContents[2648] = 8'b00000000;
        rContents[2649] = 8'b00000000;
        rContents[2650] = 8'b00000000;
        rContents[2651] = 8'b00000000;
        rContents[2652] = 8'b00000000;
        rContents[2653] = 8'b00000000;
        rContents[2654] = 8'b00000000;
        rContents[2655] = 8'b00000000;
        rContents[2656] = 8'b00000000;
        rContents[2657] = 8'b00000000;
        rContents[2658] = 8'b00000000;
        rContents[2659] = 8'b00000000;
        rContents[2660] = 8'b00000000;
        rContents[2661] = 8'b00000000;
        rContents[2662] = 8'b00000000;
        rContents[2663] = 8'b11111110;
        rContents[2664] = 8'b00000000;
        rContents[2665] = 8'b00000000;
        rContents[2666] = 8'b00000000;
        rContents[2667] = 8'b00000000;
        rContents[2668] = 8'b00000000;
        rContents[2669] = 8'b00000000;
        rContents[2670] = 8'b00000000;
        rContents[2671] = 8'b00000000;
        rContents[2672] = 8'b10000000;
        rContents[2673] = 8'b00000010;
        rContents[2674] = 8'b00000000;
        rContents[2675] = 8'b00000000;
        rContents[2676] = 8'b00000000;
        rContents[2677] = 8'b00000000;
        rContents[2678] = 8'b00000000;
        rContents[2679] = 8'b00000000;
        rContents[2680] = 8'b00000000;
        rContents[2681] = 8'b11111110;
        rContents[2682] = 8'b00000000;
        rContents[2683] = 8'b00000000;
        rContents[2684] = 8'b00000000;
        rContents[2685] = 8'b00000000;
        rContents[2686] = 8'b00000000;
        rContents[2687] = 8'b00000000;
        rContents[2688] = 8'b00000000;
        rContents[2689] = 8'b11110000;
        rContents[2690] = 8'b00001111;
        rContents[2691] = 8'b11111111;
        rContents[2692] = 8'b11111111;
        rContents[2693] = 8'b00000000;
        rContents[2694] = 8'b00000000;
        rContents[2695] = 8'b11110000;
        rContents[2696] = 8'b00001111;
        rContents[2697] = 8'b11110000;
        rContents[2698] = 8'b00001111;
        rContents[2699] = 8'b00000000;
        rContents[2700] = 8'b11111111;
        rContents[2701] = 8'b00011000;
        rContents[2702] = 8'b00000000;
        rContents[2703] = 8'b00011000;
        rContents[2704] = 8'b00000000;
        rContents[2705] = 8'b00011000;
        rContents[2706] = 8'b00011000;
        rContents[2707] = 8'b00000000;
        rContents[2708] = 8'b00011000;
        rContents[2709] = 8'b00000000;
        rContents[2710] = 8'b00011000;
        rContents[2711] = 8'b00011000;
        rContents[2712] = 8'b00100100;
        rContents[2713] = 8'b00000000;
        rContents[2714] = 8'b00100100;
        rContents[2715] = 8'b00000000;
        rContents[2716] = 8'b00100100;
        rContents[2717] = 8'b00100100;
        rContents[2718] = 8'b00000000;
        rContents[2719] = 8'b00100100;
        rContents[2720] = 8'b00100100;
        rContents[2721] = 8'b00100100;
        rContents[2722] = 8'b00000000;
        rContents[2723] = 8'b00000000;
        rContents[2724] = 8'b00000000;
        rContents[2725] = 8'b00000000;
        rContents[2726] = 8'b00000000;
        rContents[2727] = 8'b00000000;
        rContents[2728] = 8'b00000000;
        rContents[2729] = 8'b00000000;
        rContents[2730] = 8'b00000000;
        rContents[2731] = 8'b00000000;
        rContents[2732] = 8'b00000000;
        rContents[2733] = 8'b00000000;
        rContents[2734] = 8'b00000000;
        rContents[2735] = 8'b00000000;
        rContents[2736] = 8'b00000000;
        rContents[2737] = 8'b00000000;
        rContents[2738] = 8'b00000000;
        rContents[2739] = 8'b00000000;
        rContents[2740] = 8'b00000000;
        rContents[2741] = 8'b00000000;
        rContents[2742] = 8'b00000000;
        rContents[2743] = 8'b00000000;
        rContents[2744] = 8'b00000000;
        rContents[2745] = 8'b00000000;
        rContents[2746] = 8'b00000000;
        rContents[2747] = 8'b00000000;
        rContents[2748] = 8'b00000000;
        rContents[2749] = 8'b00000000;
        rContents[2750] = 8'b00000000;
        rContents[2751] = 8'b00000000;
        rContents[2752] = 8'b00000000;
        rContents[2753] = 8'b00000000;
        rContents[2754] = 8'b00000000;
        rContents[2755] = 8'b00000000;
        rContents[2756] = 8'b00000000;
        rContents[2757] = 8'b00000000;
        rContents[2758] = 8'b00000000;
        rContents[2759] = 8'b00000000;
        rContents[2760] = 8'b00000000;
        rContents[2761] = 8'b00000000;
        rContents[2762] = 8'b00000000;
        rContents[2763] = 8'b00000000;
        rContents[2764] = 8'b00000000;
        rContents[2765] = 8'b00000000;
        rContents[2766] = 8'b00000000;
        rContents[2767] = 8'b00000000;
        rContents[2768] = 8'b00000000;
        rContents[2769] = 8'b00000000;
        rContents[2770] = 8'b00000000;
        rContents[2771] = 8'b00000000;
        rContents[2772] = 8'b00000000;
        rContents[2773] = 8'b00000000;
        rContents[2774] = 8'b00000000;
        rContents[2775] = 8'b00000000;
        rContents[2776] = 8'b00000000;
        rContents[2777] = 8'b00000000;
        rContents[2778] = 8'b00000000;
        rContents[2779] = 8'b00000000;
        rContents[2780] = 8'b00000000;
        rContents[2781] = 8'b00000000;
        rContents[2782] = 8'b00000000;
        rContents[2783] = 8'b00000000;
        rContents[2784] = 8'b00000000;
        rContents[2785] = 8'b00000000;
        rContents[2786] = 8'b00000000;
        rContents[2787] = 8'b00000000;
        rContents[2788] = 8'b00000000;
        rContents[2789] = 8'b00000000;
        rContents[2790] = 8'b00000000;
        rContents[2791] = 8'b00000000;
        rContents[2792] = 8'b00000000;
        rContents[2793] = 8'b00000000;
        rContents[2794] = 8'b00000000;
        rContents[2795] = 8'b00000000;
        rContents[2796] = 8'b00000000;
        rContents[2797] = 8'b00000000;
        rContents[2798] = 8'b00000000;
        rContents[2799] = 8'b00000000;
        rContents[2800] = 8'b00000000;
        rContents[2801] = 8'b00000000;
        rContents[2802] = 8'b00000000;
        rContents[2803] = 8'b00000000;
        rContents[2804] = 8'b00000000;
        rContents[2805] = 8'b00000000;
        rContents[2806] = 8'b00000000;
        rContents[2807] = 8'b00000000;
        rContents[2808] = 8'b00000000;
        rContents[2809] = 8'b00000000;
        rContents[2810] = 8'b00000000;
        rContents[2811] = 8'b00000000;
        rContents[2812] = 8'b00000000;
        rContents[2813] = 8'b00000000;
        rContents[2814] = 8'b00000000;
        rContents[2815] = 8'b00000000;
        rContents[2816] = 8'b01010101;
        rContents[2817] = 8'b10101010;
        rContents[2818] = 8'b11111111;
        rContents[2819] = 8'b10101010;
        rContents[2820] = 8'b11111111;
        rContents[2821] = 8'b00000000;
        rContents[2822] = 8'b00000000;
        rContents[2823] = 8'b00000000;
        rContents[2824] = 8'b00000000;
        rContents[2825] = 8'b00000000;
        rContents[2826] = 8'b00000000;
        rContents[2827] = 8'b00000000;
        rContents[2828] = 8'b00000000;
        rContents[2829] = 8'b00000000;
        rContents[2830] = 8'b00000000;
        rContents[2831] = 8'b00000000;
        rContents[2832] = 8'b00000000;
        rContents[2833] = 8'b00000000;
        rContents[2834] = 8'b00000000;
        rContents[2835] = 8'b00000000;
        rContents[2836] = 8'b00000000;
        rContents[2837] = 8'b00000000;
        rContents[2838] = 8'b00000000;
        rContents[2839] = 8'b00000000;
        rContents[2840] = 8'b00000000;
        rContents[2841] = 8'b00000000;
        rContents[2842] = 8'b00000000;
        rContents[2843] = 8'b00000000;
        rContents[2844] = 8'b00000000;
        rContents[2845] = 8'b00000000;
        rContents[2846] = 8'b00000000;
        rContents[2847] = 8'b00000000;
        rContents[2848] = 8'b00000000;
        rContents[2849] = 8'b00000000;
        rContents[2850] = 8'b00000000;
        rContents[2851] = 8'b00000000;
        rContents[2852] = 8'b00000000;
        rContents[2853] = 8'b00000000;
        rContents[2854] = 8'b00000000;
        rContents[2855] = 8'b00000000;
        rContents[2856] = 8'b00000000;
        rContents[2857] = 8'b00000000;
        rContents[2858] = 8'b00000000;
        rContents[2859] = 8'b00000000;
        rContents[2860] = 8'b00000000;
        rContents[2861] = 8'b00000000;
        rContents[2862] = 8'b00000000;
        rContents[2863] = 8'b00000000;
        rContents[2864] = 8'b00000000;
        rContents[2865] = 8'b00000000;
        rContents[2866] = 8'b00000000;
        rContents[2867] = 8'b00000000;
        rContents[2868] = 8'b00000000;
        rContents[2869] = 8'b00000000;
        rContents[2870] = 8'b00000000;
        rContents[2871] = 8'b00000000;
        rContents[2872] = 8'b00000000;
        rContents[2873] = 8'b00000000;
        rContents[2874] = 8'b00000000;
        rContents[2875] = 8'b00000000;
        rContents[2876] = 8'b00000000;
        rContents[2877] = 8'b00000000;
        rContents[2878] = 8'b00000000;
        rContents[2879] = 8'b00000000;
        rContents[2880] = 8'b00000000;
        rContents[2881] = 8'b00000000;
        rContents[2882] = 8'b00000000;
        rContents[2883] = 8'b00000000;
        rContents[2884] = 8'b00000000;
        rContents[2885] = 8'b00000000;
        rContents[2886] = 8'b00000000;
        rContents[2887] = 8'b00000000;
        rContents[2888] = 8'b00000000;
        rContents[2889] = 8'b00000000;
        rContents[2890] = 8'b00000000;
        rContents[2891] = 8'b00000000;
        rContents[2892] = 8'b00000000;
        rContents[2893] = 8'b00000000;
        rContents[2894] = 8'b00000000;
        rContents[2895] = 8'b00000000;
        rContents[2896] = 8'b00000000;
        rContents[2897] = 8'b00000000;
        rContents[2898] = 8'b00000000;
        rContents[2899] = 8'b00000000;
        rContents[2900] = 8'b00000000;
        rContents[2901] = 8'b00000000;
        rContents[2902] = 8'b00000000;
        rContents[2903] = 8'b00000000;
        rContents[2904] = 8'b00000000;
        rContents[2905] = 8'b00000000;
        rContents[2906] = 8'b00000000;
        rContents[2907] = 8'b00000000;
        rContents[2908] = 8'b00000000;
        rContents[2909] = 8'b00000000;
        rContents[2910] = 8'b00000000;
        rContents[2911] = 8'b00000000;
        rContents[2912] = 8'b00000000;
        rContents[2913] = 8'b00000000;
        rContents[2914] = 8'b00000000;
        rContents[2915] = 8'b00000000;
        rContents[2916] = 8'b00000000;
        rContents[2917] = 8'b00000000;
        rContents[2918] = 8'b00000000;
        rContents[2919] = 8'b00000000;
        rContents[2920] = 8'b00000000;
        rContents[2921] = 8'b00000000;
        rContents[2922] = 8'b00000000;
        rContents[2923] = 8'b00000000;
        rContents[2924] = 8'b00000000;
        rContents[2925] = 8'b00000000;
        rContents[2926] = 8'b00000000;
        rContents[2927] = 8'b00000000;
        rContents[2928] = 8'b00000000;
        rContents[2929] = 8'b00000000;
        rContents[2930] = 8'b00000000;
        rContents[2931] = 8'b00000000;
        rContents[2932] = 8'b00000000;
        rContents[2933] = 8'b00000000;
        rContents[2934] = 8'b00000000;
        rContents[2935] = 8'b00000000;
        rContents[2936] = 8'b00000000;
        rContents[2937] = 8'b00000000;
        rContents[2938] = 8'b00000000;
        rContents[2939] = 8'b00000000;
        rContents[2940] = 8'b00000000;
        rContents[2941] = 8'b00000000;
        rContents[2942] = 8'b00000000;
        rContents[2943] = 8'b00000000;
        rContents[2944] = 8'b00000000;
        rContents[2945] = 8'b11110000;
        rContents[2946] = 8'b00001111;
        rContents[2947] = 8'b11111111;
        rContents[2948] = 8'b11111111;
        rContents[2949] = 8'b00000000;
        rContents[2950] = 8'b00000000;
        rContents[2951] = 8'b11110000;
        rContents[2952] = 8'b00001111;
        rContents[2953] = 8'b11110000;
        rContents[2954] = 8'b00001111;
        rContents[2955] = 8'b00000000;
        rContents[2956] = 8'b11111111;
        rContents[2957] = 8'b00011000;
        rContents[2958] = 8'b00000000;
        rContents[2959] = 8'b00011000;
        rContents[2960] = 8'b00000000;
        rContents[2961] = 8'b00011000;
        rContents[2962] = 8'b00011000;
        rContents[2963] = 8'b00000000;
        rContents[2964] = 8'b00011000;
        rContents[2965] = 8'b00000000;
        rContents[2966] = 8'b00011000;
        rContents[2967] = 8'b00011000;
        rContents[2968] = 8'b00100100;
        rContents[2969] = 8'b00000000;
        rContents[2970] = 8'b00100100;
        rContents[2971] = 8'b00000000;
        rContents[2972] = 8'b00100100;
        rContents[2973] = 8'b00100100;
        rContents[2974] = 8'b00000000;
        rContents[2975] = 8'b00100100;
        rContents[2976] = 8'b00100100;
        rContents[2977] = 8'b00100100;
        rContents[2978] = 8'b00000000;
        rContents[2979] = 8'b00000000;
        rContents[2980] = 8'b00000000;
        rContents[2981] = 8'b00000000;
        rContents[2982] = 8'b00000000;
        rContents[2983] = 8'b00000000;
        rContents[2984] = 8'b00000000;
        rContents[2985] = 8'b00000000;
        rContents[2986] = 8'b00000000;
        rContents[2987] = 8'b00000000;
        rContents[2988] = 8'b00000000;
        rContents[2989] = 8'b00000000;
        rContents[2990] = 8'b00000000;
        rContents[2991] = 8'b00000000;
        rContents[2992] = 8'b00000000;
        rContents[2993] = 8'b00000000;
        rContents[2994] = 8'b00000000;
        rContents[2995] = 8'b00000000;
        rContents[2996] = 8'b00000000;
        rContents[2997] = 8'b00000000;
        rContents[2998] = 8'b00000000;
        rContents[2999] = 8'b00000000;
        rContents[3000] = 8'b00000000;
        rContents[3001] = 8'b00000000;
        rContents[3002] = 8'b00000000;
        rContents[3003] = 8'b00000000;
        rContents[3004] = 8'b00000000;
        rContents[3005] = 8'b00000000;
        rContents[3006] = 8'b00000000;
        rContents[3007] = 8'b00000000;
        rContents[3008] = 8'b00000000;
        rContents[3009] = 8'b00000000;
        rContents[3010] = 8'b00000000;
        rContents[3011] = 8'b00000000;
        rContents[3012] = 8'b00000000;
        rContents[3013] = 8'b00000000;
        rContents[3014] = 8'b00000000;
        rContents[3015] = 8'b00000000;
        rContents[3016] = 8'b00000000;
        rContents[3017] = 8'b00000000;
        rContents[3018] = 8'b00000000;
        rContents[3019] = 8'b00000000;
        rContents[3020] = 8'b00000000;
        rContents[3021] = 8'b00000000;
        rContents[3022] = 8'b00000000;
        rContents[3023] = 8'b00000000;
        rContents[3024] = 8'b00000000;
        rContents[3025] = 8'b00000000;
        rContents[3026] = 8'b00000000;
        rContents[3027] = 8'b00000000;
        rContents[3028] = 8'b00000000;
        rContents[3029] = 8'b00000000;
        rContents[3030] = 8'b00000000;
        rContents[3031] = 8'b00000000;
        rContents[3032] = 8'b00000000;
        rContents[3033] = 8'b00000000;
        rContents[3034] = 8'b00000000;
        rContents[3035] = 8'b00000000;
        rContents[3036] = 8'b00000000;
        rContents[3037] = 8'b00000000;
        rContents[3038] = 8'b00000000;
        rContents[3039] = 8'b00000000;
        rContents[3040] = 8'b00000000;
        rContents[3041] = 8'b00000000;
        rContents[3042] = 8'b00000000;
        rContents[3043] = 8'b00000000;
        rContents[3044] = 8'b00000000;
        rContents[3045] = 8'b00000000;
        rContents[3046] = 8'b00000000;
        rContents[3047] = 8'b00000000;
        rContents[3048] = 8'b00000000;
        rContents[3049] = 8'b00000000;
        rContents[3050] = 8'b00000000;
        rContents[3051] = 8'b00000000;
        rContents[3052] = 8'b00000000;
        rContents[3053] = 8'b00000000;
        rContents[3054] = 8'b00000000;
        rContents[3055] = 8'b00000000;
        rContents[3056] = 8'b00000000;
        rContents[3057] = 8'b00000000;
        rContents[3058] = 8'b00000000;
        rContents[3059] = 8'b00000000;
        rContents[3060] = 8'b00000000;
        rContents[3061] = 8'b00000000;
        rContents[3062] = 8'b00000000;
        rContents[3063] = 8'b00000000;
        rContents[3064] = 8'b00000000;
        rContents[3065] = 8'b00000000;
        rContents[3066] = 8'b00000000;
        rContents[3067] = 8'b00000000;
        rContents[3068] = 8'b00000000;
        rContents[3069] = 8'b00000000;
        rContents[3070] = 8'b00000000;
        rContents[3071] = 8'b00000000;
    end
    
endmodule
