module epRISC_embeddedROM(iClk, iAddr, oData, iEnable);

    input iClk, iEnable;
    input [11:0] iAddr;
    output wire [31:0] oData;
    
    reg [31:0] rDataOut, rContents[0:4095];
    
    assign oData = (iEnable) ? rDataOut : 32'bz;
    
    always @(posedge iClk) begin
        rDataOut = rContents[iAddr];
    end
    
    initial begin
rContents[0] = 32'h21001100;
rContents[1] = 32'h23000000;
rContents[2] = 32'hD00000FF;
rContents[3] = 32'h24007FFF;
rContents[4] = 32'h61400000;
rContents[5] = 32'h24000000;
rContents[6] = 32'h61400000;
rContents[7] = 32'hD0000107;
rContents[8] = 32'h41400000;
rContents[9] = 32'h41400000;
rContents[10] = 32'h240000FF;
rContents[11] = 32'h61400000;
rContents[12] = 32'hD0000364;
rContents[13] = 32'h41400000;
rContents[14] = 32'h2400004B;
rContents[15] = 32'h61400000;
rContents[16] = 32'hD00001FA;
rContents[17] = 32'h41400000;
rContents[18] = 32'h240000CD;
rContents[19] = 32'h61400000;
rContents[20] = 32'hD00001F6;
rContents[21] = 32'h41400000;
rContents[22] = 32'h240000EF;
rContents[23] = 32'h61400000;
rContents[24] = 32'hD00001F2;
rContents[25] = 32'h41400000;
rContents[26] = 32'h24000041;
rContents[27] = 32'h61400000;
rContents[28] = 32'hD0000181;
rContents[29] = 32'h41400000;
rContents[30] = 32'h2400005C;
rContents[31] = 32'h61400000;
rContents[32] = 32'hD00001EA;
rContents[33] = 32'h41400000;
rContents[34] = 32'hD00001FE;
rContents[35] = 32'h2400007B;
rContents[36] = 32'h18E0F0FF;
rContents[37] = 32'h81000002;
rContents[38] = 32'h24000072;
rContents[39] = 32'h61400000;
rContents[40] = 32'hD00001E2;
rContents[41] = 32'h41400000;
rContents[42] = 32'h24003000;
rContents[43] = 32'h61400000;
rContents[44] = 32'h24000000;
rContents[45] = 32'h61400000;
rContents[46] = 32'hD00002C2;
rContents[47] = 32'h41400000;
rContents[48] = 32'h41400000;
rContents[49] = 32'h240000FB;
rContents[50] = 32'h61400000;
rContents[51] = 32'hD00001D7;
rContents[52] = 32'h41400000;
rContents[53] = 32'h80000427;
rContents[54] = 32'h43F01FF0;
rContents[55] = 32'h61F00000;
rContents[56] = 32'hD0000165;
rContents[57] = 32'h63F01FF1;
rContents[58] = 32'h41F00000;
rContents[59] = 32'hF0000000;
rContents[60] = 32'hD0000183;
rContents[61] = 32'h63F01FF1;
rContents[62] = 32'hF0000000;
rContents[63] = 32'h43F01FF2;
rContents[64] = 32'h61F00000;
rContents[65] = 32'h43F01FF3;
rContents[66] = 32'h61F00000;
rContents[67] = 32'hD0000278;
rContents[68] = 32'h63F01FF4;
rContents[69] = 32'h41F00000;
rContents[70] = 32'h41F00000;
rContents[71] = 32'hF0000000;
rContents[72] = 32'hD00001D8;
rContents[73] = 32'h63F01FF5;
rContents[74] = 32'hF0000000;
rContents[75] = 32'h65705249;
rContents[76] = 32'h53432042;
rContents[77] = 32'h6F6F746C;
rContents[78] = 32'h6F616465;
rContents[79] = 32'h72207633;
rContents[80] = 32'h2E320A0D;
rContents[81] = 32'h636F7079;
rContents[82] = 32'h72696768;
rContents[83] = 32'h74203230;
rContents[84] = 32'h31352D32;
rContents[85] = 32'h30313720;
rContents[86] = 32'h50726F70;
rContents[87] = 32'h6F727469;
rContents[88] = 32'h6F6E616C;
rContents[89] = 32'h204C6162;
rContents[90] = 32'h730A0D0A;
rContents[91] = 32'h0D000000;
rContents[92] = 32'h41747465;
rContents[93] = 32'h6D707469;
rContents[94] = 32'h6E672074;
rContents[95] = 32'h6F206D6F;
rContents[96] = 32'h756E7420;
rContents[97] = 32'h53442063;
rContents[98] = 32'h61726420;
rContents[99] = 32'h696E2073;
rContents[100] = 32'h6C6F7420;
rContents[101] = 32'h412E2E2E;
rContents[102] = 32'h0A0D0000;
rContents[103] = 32'h41747465;
rContents[104] = 32'h6D707469;
rContents[105] = 32'h6E672074;
rContents[106] = 32'h6F206D6F;
rContents[107] = 32'h756E7420;
rContents[108] = 32'h53442063;
rContents[109] = 32'h61726420;
rContents[110] = 32'h696E2073;
rContents[111] = 32'h6C6F7420;
rContents[112] = 32'h422E2E2E;
rContents[113] = 32'h0A0D0000;
rContents[114] = 32'h20205344;
rContents[115] = 32'h20636172;
rContents[116] = 32'h64206D6F;
rContents[117] = 32'h756E7465;
rContents[118] = 32'h64207375;
rContents[119] = 32'h63636573;
rContents[120] = 32'h7366756C;
rContents[121] = 32'h6C792E0A;
rContents[122] = 32'h0D0A0D00;
rContents[123] = 32'h20204572;
rContents[124] = 32'h726F7220;
rContents[125] = 32'h6D6F756E;
rContents[126] = 32'h74696E67;
rContents[127] = 32'h20534420;
rContents[128] = 32'h63617264;
rContents[129] = 32'h2E0A0D0A;
rContents[130] = 32'h0D000000;
rContents[131] = 32'h46657463;
rContents[132] = 32'h68696E67;
rContents[133] = 32'h20646973;
rContents[134] = 32'h6B20696E;
rContents[135] = 32'h666F2E2E;
rContents[136] = 32'h2E0A0D00;
rContents[137] = 32'h20204469;
rContents[138] = 32'h736B2061;
rContents[139] = 32'h70706561;
rContents[140] = 32'h72732074;
rContents[141] = 32'h6F206265;
rContents[142] = 32'h20636F72;
rContents[143] = 32'h72757074;
rContents[144] = 32'h2E0A0D0A;
rContents[145] = 32'h0D000000;
rContents[146] = 32'h2020466F;
rContents[147] = 32'h756E6420;
rContents[148] = 32'h6469736B;
rContents[149] = 32'h20270000;
rContents[150] = 32'h27206174;
rContents[151] = 32'h20626C6F;
rContents[152] = 32'h636B2030;
rContents[153] = 32'h2E0A0D00;
rContents[154] = 32'h20204469;
rContents[155] = 32'h736B2061;
rContents[156] = 32'h70706561;
rContents[157] = 32'h72732074;
rContents[158] = 32'h6F206265;
rContents[159] = 32'h20656D70;
rContents[160] = 32'h74792E0A;
rContents[161] = 32'h0D0A0D00;
rContents[162] = 32'h2020466F;
rContents[163] = 32'h756E6420;
rContents[164] = 32'h00000000;
rContents[165] = 32'h20656E74;
rContents[166] = 32'h72696573;
rContents[167] = 32'h206F6E20;
rContents[168] = 32'h6469736B;
rContents[169] = 32'h2E0A0D0A;
rContents[170] = 32'h0D000000;
rContents[171] = 32'h41766169;
rContents[172] = 32'h6C61626C;
rContents[173] = 32'h6520656E;
rContents[174] = 32'h74726965;
rContents[175] = 32'h733A0A0D;
rContents[176] = 32'h00000000;
rContents[177] = 32'h2020456E;
rContents[178] = 32'h74727920;
rContents[179] = 32'h27000000;
rContents[180] = 32'h273A2073;
rContents[181] = 32'h74617274;
rContents[182] = 32'h20000000;
rContents[183] = 32'h2C206C65;
rContents[184] = 32'h6E677468;
rContents[185] = 32'h20000000;
rContents[186] = 32'h2C206C6F;
rContents[187] = 32'h6164200A;
rContents[188] = 32'h0D000000;
rContents[189] = 32'h53656C65;
rContents[190] = 32'h63742061;
rContents[191] = 32'h6E20656E;
rContents[192] = 32'h74727920;
rContents[193] = 32'h746F2065;
rContents[194] = 32'h78656375;
rContents[195] = 32'h74652C20;
rContents[196] = 32'h6F722074;
rContents[197] = 32'h79706520;
rContents[198] = 32'h276D2720;
rContents[199] = 32'h746F2065;
rContents[200] = 32'h6E746572;
rContents[201] = 32'h20746865;
rContents[202] = 32'h206D6F6E;
rContents[203] = 32'h69746F72;
rContents[204] = 32'h3A000000;
rContents[205] = 32'h53746172;
rContents[206] = 32'h74696E67;
rContents[207] = 32'h20504F53;
rContents[208] = 32'h54732E2E;
rContents[209] = 32'h2E0A0D00;
rContents[210] = 32'h20204D65;
rContents[211] = 32'h6D6F7279;
rContents[212] = 32'h20202020;
rContents[213] = 32'h20202020;
rContents[214] = 32'h20200000;
rContents[215] = 32'h20205541;
rContents[216] = 32'h52542020;
rContents[217] = 32'h20202020;
rContents[218] = 32'h20202020;
rContents[219] = 32'h20200000;
rContents[220] = 32'h20205350;
rContents[221] = 32'h49202020;
rContents[222] = 32'h20202020;
rContents[223] = 32'h20202020;
rContents[224] = 32'h20200000;
rContents[225] = 32'h20207379;
rContents[226] = 32'h73582042;
rContents[227] = 32'h75732020;
rContents[228] = 32'h20202020;
rContents[229] = 32'h20200000;
rContents[230] = 32'h2020492F;
rContents[231] = 32'h4F20436F;
rContents[232] = 32'h6E74726F;
rContents[233] = 32'h6C6C6572;
rContents[234] = 32'h20200000;
rContents[235] = 32'h4F4B0A0D;
rContents[236] = 32'h00000000;
rContents[237] = 32'h4641494C;
rContents[238] = 32'h0A0D0000;
rContents[239] = 32'h504F5354;
rContents[240] = 32'h20737563;
rContents[241] = 32'h63657373;
rContents[242] = 32'h66756C2E;
rContents[243] = 32'h0A0D0A0D;
rContents[244] = 32'h00000000;
rContents[245] = 32'h504F5354;
rContents[246] = 32'h20756E73;
rContents[247] = 32'h75636365;
rContents[248] = 32'h73736675;
rContents[249] = 32'h6C2E0A0D;
rContents[250] = 32'h0A0D0000;
rContents[251] = 32'h456E7465;
rContents[252] = 32'h72696E67;
rContents[253] = 32'h206D6F6E;
rContents[254] = 32'h69746F72;
rContents[255] = 32'h2E2E2E0A;
rContents[256] = 32'h0D0A0D00;
rContents[257] = 32'h61C00000;
rContents[258] = 32'h2C002000;
rContents[259] = 32'h2F010001;
rContents[260] = 32'h6CF00000;
rContents[261] = 32'h04000000;
rContents[262] = 32'h04000000;
rContents[263] = 32'h04000000;
rContents[264] = 32'h04000000;
rContents[265] = 32'h4CF00000;
rContents[266] = 32'h18F0F001;
rContents[267] = 32'h820FFFFE;
rContents[268] = 32'h41C00000;
rContents[269] = 32'hF0000000;
rContents[270] = 32'h61E00000;
rContents[271] = 32'h61D00000;
rContents[272] = 32'h61C00000;
rContents[273] = 32'h18111004;
rContents[274] = 32'h2C002000;
rContents[275] = 32'h41D00000;
rContents[276] = 32'h41E00000;
rContents[277] = 32'h18011006;
rContents[278] = 32'h2F600008;
rContents[279] = 32'h103FFE00;
rContents[280] = 32'h186FF010;
rContents[281] = 32'h103FFD00;
rContents[282] = 32'h6CF00001;
rContents[283] = 32'h2F010005;
rContents[284] = 32'h6CF00000;
rContents[285] = 32'h4CF00000;
rContents[286] = 32'h18F0F001;
rContents[287] = 32'h820FFFFE;
rContents[288] = 32'h4CF00002;
rContents[289] = 32'h41C00000;
rContents[290] = 32'h41D00000;
rContents[291] = 32'h41E00000;
rContents[292] = 32'hF0000000;
rContents[293] = 32'h61E00000;
rContents[294] = 32'h61C00000;
rContents[295] = 32'h18111003;
rContents[296] = 32'h2C002000;
rContents[297] = 32'h41E00000;
rContents[298] = 32'h18011004;
rContents[299] = 32'h2F600000;
rContents[300] = 32'h103FFE00;
rContents[301] = 32'h186FF010;
rContents[302] = 32'h6CF00001;
rContents[303] = 32'h2F010005;
rContents[304] = 32'h6CF00000;
rContents[305] = 32'h4CF00000;
rContents[306] = 32'h18F0F001;
rContents[307] = 32'h820FFFFE;
rContents[308] = 32'h2F600000;
rContents[309] = 32'h103FFE00;
rContents[310] = 32'h186FF010;
rContents[311] = 32'h6CF00001;
rContents[312] = 32'h2F010005;
rContents[313] = 32'h6CF00000;
rContents[314] = 32'h4CF00000;
rContents[315] = 32'h18F0F001;
rContents[316] = 32'h820FFFFE;
rContents[317] = 32'h4CF00002;
rContents[318] = 32'h41C00000;
rContents[319] = 32'h41E00000;
rContents[320] = 32'hF0000000;
rContents[321] = 32'h61D00000;
rContents[322] = 32'h61C00000;
rContents[323] = 32'h18111003;
rContents[324] = 32'h2C002000;
rContents[325] = 32'h41D00000;
rContents[326] = 32'h18011004;
rContents[327] = 32'h2F000011;
rContents[328] = 32'h61F00000;
rContents[329] = 32'h61D00000;
rContents[330] = 32'hD00FFFC4;
rContents[331] = 32'h41D00000;
rContents[332] = 32'h41F00000;
rContents[333] = 32'h2F000010;
rContents[334] = 32'h61F00000;
rContents[335] = 32'h2F000080;
rContents[336] = 32'h61F00000;
rContents[337] = 32'hD00FFFBD;
rContents[338] = 32'h41D00000;
rContents[339] = 32'h41F00000;
rContents[340] = 32'h2F000010;
rContents[341] = 32'h61F00000;
rContents[342] = 32'hD00FFFCF;
rContents[343] = 32'h18F0F080;
rContents[344] = 32'h820FFFFE;
rContents[345] = 32'h41F00000;
rContents[346] = 32'h41C00000;
rContents[347] = 32'h41D00000;
rContents[348] = 32'hF0000000;
rContents[349] = 32'h61C00000;
rContents[350] = 32'h2C002000;
rContents[351] = 32'h2F808010;
rContents[352] = 32'h3F000020;
rContents[353] = 32'h6CF00001;
rContents[354] = 32'h2F010005;
rContents[355] = 32'h6CF00000;
rContents[356] = 32'h4CF00000;
rContents[357] = 32'h18F0F001;
rContents[358] = 32'h820FFFFE;
rContents[359] = 32'h2F800010;
rContents[360] = 32'h6CF00001;
rContents[361] = 32'h2F010005;
rContents[362] = 32'h6CF00000;
rContents[363] = 32'h4CF00000;
rContents[364] = 32'h18F0F001;
rContents[365] = 32'h820FFFFE;
rContents[366] = 32'h2F800010;
rContents[367] = 32'h6CF00001;
rContents[368] = 32'h2F010005;
rContents[369] = 32'h6CF00000;
rContents[370] = 32'h4CF00000;
rContents[371] = 32'h18F0F001;
rContents[372] = 32'h820FFFFE;
rContents[373] = 32'h4CF00002;
rContents[374] = 32'h18F0F020;
rContents[375] = 32'h820FFFF7;
rContents[376] = 32'h2F800012;
rContents[377] = 32'h6CF00001;
rContents[378] = 32'h2F010005;
rContents[379] = 32'h6CF00000;
rContents[380] = 32'h4CF00000;
rContents[381] = 32'h18F0F001;
rContents[382] = 32'h820FFFFE;
rContents[383] = 32'h2F800012;
rContents[384] = 32'h6CF00001;
rContents[385] = 32'h2F010005;
rContents[386] = 32'h6CF00000;
rContents[387] = 32'h4CF00000;
rContents[388] = 32'h18F0F001;
rContents[389] = 32'h820FFFFE;
rContents[390] = 32'h4CF00002;
rContents[391] = 32'h41C00000;
rContents[392] = 32'hF0000000;
rContents[393] = 32'h61C00000;
rContents[394] = 32'h61D00000;
rContents[395] = 32'h18111003;
rContents[396] = 32'h41C00000;
rContents[397] = 32'h18011004;
rContents[398] = 32'h2D000020;
rContents[399] = 32'h61D00000;
rContents[400] = 32'hD00FFF95;
rContents[401] = 32'h41D00000;
rContents[402] = 32'h18BFF078;
rContents[403] = 32'h186CC003;
rContents[404] = 32'h103CCF00;
rContents[405] = 32'h61D00000;
rContents[406] = 32'h61C00000;
rContents[407] = 32'hD00FFF77;
rContents[408] = 32'h41C00000;
rContents[409] = 32'h41D00000;
rContents[410] = 32'h41D00000;
rContents[411] = 32'h41C00000;
rContents[412] = 32'hF0000000;
rContents[413] = 32'h61C00000;
rContents[414] = 32'h61D00000;
rContents[415] = 32'h18111003;
rContents[416] = 32'h41C00000;
rContents[417] = 32'h18011004;
rContents[418] = 32'h2D000021;
rContents[419] = 32'h61D00000;
rContents[420] = 32'h61C00000;
rContents[421] = 32'hD00FFF69;
rContents[422] = 32'h41C00000;
rContents[423] = 32'h41D00000;
rContents[424] = 32'h2D000020;
rContents[425] = 32'h61D00000;
rContents[426] = 32'hD00FFF7B;
rContents[427] = 32'h41D00000;
rContents[428] = 32'h183FF080;
rContents[429] = 32'h61D00000;
rContents[430] = 32'h61F00000;
rContents[431] = 32'hD00FFF5F;
rContents[432] = 32'h41F00000;
rContents[433] = 32'h41D00000;
rContents[434] = 32'h2D000020;
rContents[435] = 32'h61D00000;
rContents[436] = 32'hD00FFF71;
rContents[437] = 32'h18F0F080;
rContents[438] = 32'h820FFFFE;
rContents[439] = 32'h41D00000;
rContents[440] = 32'h2D000022;
rContents[441] = 32'h61D00000;
rContents[442] = 32'hD00FFF6B;
rContents[443] = 32'h41D00000;
rContents[444] = 32'h41D00000;
rContents[445] = 32'h41C00000;
rContents[446] = 32'hF0000000;
rContents[447] = 32'h61D00000;
rContents[448] = 32'h2D000021;
rContents[449] = 32'h61D00000;
rContents[450] = 32'h2D0000FF;
rContents[451] = 32'h61D00000;
rContents[452] = 32'hD00FFF4A;
rContents[453] = 32'h41D00000;
rContents[454] = 32'h41D00000;
rContents[455] = 32'h2D000020;
rContents[456] = 32'h61D00000;
rContents[457] = 32'hD00FFF5C;
rContents[458] = 32'h41D00000;
rContents[459] = 32'h183FF080;
rContents[460] = 32'h61D00000;
rContents[461] = 32'h61F00000;
rContents[462] = 32'hD00FFF40;
rContents[463] = 32'h41F00000;
rContents[464] = 32'h41D00000;
rContents[465] = 32'h2D000020;
rContents[466] = 32'h61D00000;
rContents[467] = 32'hD00FFF52;
rContents[468] = 32'h18F0F080;
rContents[469] = 32'h820FFFFE;
rContents[470] = 32'h41D00000;
rContents[471] = 32'h2D000022;
rContents[472] = 32'h61D00000;
rContents[473] = 32'hD00FFF4C;
rContents[474] = 32'h41D00000;
rContents[475] = 32'h41D00000;
rContents[476] = 32'hF0000000;
rContents[477] = 32'h61C00000;
rContents[478] = 32'h61D00000;
rContents[479] = 32'h61E00000;
rContents[480] = 32'h18111004;
rContents[481] = 32'h41C00000;
rContents[482] = 32'h2E000008;
rContents[483] = 32'h18011005;
rContents[484] = 32'h182DCCF0;
rContents[485] = 32'h186CC004;
rContents[486] = 32'h188DD01C;
rContents[487] = 32'h180DD030;
rContents[488] = 32'h18E0D03A;
rContents[489] = 32'h84000003;
rContents[490] = 32'h18B22008;
rContents[491] = 32'h180DD007;
rContents[492] = 32'h61D00000;
rContents[493] = 32'hD00FFF54;
rContents[494] = 32'h41D00000;
rContents[495] = 32'h181EE001;
rContents[496] = 32'h18E0E000;
rContents[497] = 32'h820FFFF3;
rContents[498] = 32'h41E00000;
rContents[499] = 32'h41D00000;
rContents[500] = 32'h41C00000;
rContents[501] = 32'hF0000000;
rContents[502] = 32'h61C00000;
rContents[503] = 32'h61D00000;
rContents[504] = 32'h61E00000;
rContents[505] = 32'h18111004;
rContents[506] = 32'h41D00000;
rContents[507] = 32'h41C00000;
rContents[508] = 32'h18011006;
rContents[509] = 32'h08ED0000;
rContents[510] = 32'h187DD002;
rContents[511] = 32'h100CCD00;
rContents[512] = 32'h4CF00000;
rContents[513] = 32'h2D000003;
rContents[514] = 32'h182EE003;
rContents[515] = 32'h101EDE00;
rContents[516] = 32'h186EE003;
rContents[517] = 32'h10DFFEFF;
rContents[518] = 32'h41E00000;
rContents[519] = 32'h41D00000;
rContents[520] = 32'h41C00000;
rContents[521] = 32'hF0000000;
rContents[522] = 32'h61C00000;
rContents[523] = 32'h61D00000;
rContents[524] = 32'h18111003;
rContents[525] = 32'h2D000000;
rContents[526] = 32'h41C00000;
rContents[527] = 32'h18011004;
rContents[528] = 32'h61C00000;
rContents[529] = 32'h61D00000;
rContents[530] = 32'hD00FFFE4;
rContents[531] = 32'h41D00000;
rContents[532] = 32'h18E0F000;
rContents[533] = 32'h81000007;
rContents[534] = 32'h61F00000;
rContents[535] = 32'hD00FFF2A;
rContents[536] = 32'hD00001AB;
rContents[537] = 32'h41F00000;
rContents[538] = 32'h180DD001;
rContents[539] = 32'h800FFFF6;
rContents[540] = 32'h41C00000;
rContents[541] = 32'h41D00000;
rContents[542] = 32'h41C00000;
rContents[543] = 32'hF0000000;
rContents[544] = 32'h61C00000;
rContents[545] = 32'h61D00000;
rContents[546] = 32'h61E00000;
rContents[547] = 32'h2C000000;
rContents[548] = 32'h61C00000;
rContents[549] = 32'hD00FFF64;
rContents[550] = 32'h41C00000;
rContents[551] = 32'h2C00000B;
rContents[552] = 32'hD00FFF97;
rContents[553] = 32'h181CC001;
rContents[554] = 32'h18E0C000;
rContents[555] = 32'h820FFFFD;
rContents[556] = 32'h2C000001;
rContents[557] = 32'h61C00000;
rContents[558] = 32'hD00FFF5B;
rContents[559] = 32'h41C00000;
rContents[560] = 32'h2C000000;
rContents[561] = 32'h61C00000;
rContents[562] = 32'h2C000000;
rContents[563] = 32'h61C00000;
rContents[564] = 32'h2D000001;
rContents[565] = 32'h186DD000;
rContents[566] = 32'h2E000000;
rContents[567] = 32'hD0000084;
rContents[568] = 32'h10E0FD00;
rContents[569] = 32'h81000005;
rContents[570] = 32'h180EE001;
rContents[571] = 32'h18E0E402;
rContents[572] = 32'h8100006E;
rContents[573] = 32'h800FFFFA;
rContents[574] = 32'h41C00000;
rContents[575] = 32'h41C00000;
rContents[576] = 32'h2C000008;
rContents[577] = 32'h61C00000;
rContents[578] = 32'h2C0001AA;
rContents[579] = 32'h61C00000;
rContents[580] = 32'hD0000077;
rContents[581] = 32'h41C00000;
rContents[582] = 32'h41C00000;
rContents[583] = 32'h2D000001;
rContents[584] = 32'h186DD002;
rContents[585] = 32'h10F0FD00;
rContents[586] = 32'h8200000C;
rContents[587] = 32'hD00FFF74;
rContents[588] = 32'hD00FFF73;
rContents[589] = 32'hD00FFF72;
rContents[590] = 32'h18F0F001;
rContents[591] = 32'h8100005D;
rContents[592] = 32'hD00FFF6F;
rContents[593] = 32'h18E0F0AA;
rContents[594] = 32'h8200005A;
rContents[595] = 32'h2E000001;
rContents[596] = 32'h186EE001;
rContents[597] = 32'h80000014;
rContents[598] = 32'h2C000037;
rContents[599] = 32'h61C00000;
rContents[600] = 32'h2C000000;
rContents[601] = 32'h61C00000;
rContents[602] = 32'hD0000061;
rContents[603] = 32'h41C00000;
rContents[604] = 32'h41C00000;
rContents[605] = 32'h2C000029;
rContents[606] = 32'h61C00000;
rContents[607] = 32'h2C000000;
rContents[608] = 32'h61C00000;
rContents[609] = 32'hD000005A;
rContents[610] = 32'h41C00000;
rContents[611] = 32'h41C00000;
rContents[612] = 32'h2E000000;
rContents[613] = 32'h10E0FD00;
rContents[614] = 32'h82000003;
rContents[615] = 32'h2E000001;
rContents[616] = 32'h186EE000;
rContents[617] = 32'h2D000000;
rContents[618] = 32'h18F0E003;
rContents[619] = 32'h81000013;
rContents[620] = 32'h2C000037;
rContents[621] = 32'h61C00000;
rContents[622] = 32'h2C000000;
rContents[623] = 32'h61C00000;
rContents[624] = 32'hD000004B;
rContents[625] = 32'h41C00000;
rContents[626] = 32'h41C00000;
rContents[627] = 32'h2C000029;
rContents[628] = 32'h61C00000;
rContents[629] = 32'h2C000000;
rContents[630] = 32'h18F0E002;
rContents[631] = 32'h81000002;
rContents[632] = 32'h2C804000;
rContents[633] = 32'h61C00000;
rContents[634] = 32'hD0000041;
rContents[635] = 32'h41C00000;
rContents[636] = 32'h41C00000;
rContents[637] = 32'h80000008;
rContents[638] = 32'h2C000029;
rContents[639] = 32'h61C00000;
rContents[640] = 32'h2C000000;
rContents[641] = 32'h61C00000;
rContents[642] = 32'hD0000039;
rContents[643] = 32'h41C00000;
rContents[644] = 32'h41C00000;
rContents[645] = 32'h18F0F001;
rContents[646] = 32'h81000005;
rContents[647] = 32'h180DD001;
rContents[648] = 32'h18E0D480;
rContents[649] = 32'h81000023;
rContents[650] = 32'h800FFFE0;
rContents[651] = 32'h18F0E002;
rContents[652] = 32'h81000013;
rContents[653] = 32'h2C00003A;
rContents[654] = 32'h61C00000;
rContents[655] = 32'h2C000000;
rContents[656] = 32'h61C00000;
rContents[657] = 32'hD000002A;
rContents[658] = 32'h41C00000;
rContents[659] = 32'h41C00000;
rContents[660] = 32'h18E0F000;
rContents[661] = 32'h82000017;
rContents[662] = 32'hD00FFF29;
rContents[663] = 32'h18F0F040;
rContents[664] = 32'h81000004;
rContents[665] = 32'h2C000001;
rContents[666] = 32'h186CC002;
rContents[667] = 32'h103EEC00;
rContents[668] = 32'hD00FFF23;
rContents[669] = 32'hD00FFF22;
rContents[670] = 32'hD00FFF21;
rContents[671] = 32'h2C000010;
rContents[672] = 32'h61C00000;
rContents[673] = 32'h2C000200;
rContents[674] = 32'h61C00000;
rContents[675] = 32'hD0000018;
rContents[676] = 32'h41C00000;
rContents[677] = 32'h41C00000;
rContents[678] = 32'h18E0F000;
rContents[679] = 32'h82000005;
rContents[680] = 32'h8000000A;
rContents[681] = 32'hD000018D;
rContents[682] = 32'h41C00000;
rContents[683] = 32'h41C00000;
rContents[684] = 32'h2C000000;
rContents[685] = 32'h61C00000;
rContents[686] = 32'hD00FFEDB;
rContents[687] = 32'h41C00000;
rContents[688] = 32'h2F0000FF;
rContents[689] = 32'h80000006;
rContents[690] = 32'h2C000000;
rContents[691] = 32'h61C00000;
rContents[692] = 32'hD00FFED5;
rContents[693] = 32'h41C00000;
rContents[694] = 32'h08FE0000;
rContents[695] = 32'h41E00000;
rContents[696] = 32'h41D00000;
rContents[697] = 32'h41C00000;
rContents[698] = 32'hF0000000;
rContents[699] = 32'h61C00000;
rContents[700] = 32'h61D00000;
rContents[701] = 32'h18111003;
rContents[702] = 32'h41D00000;
rContents[703] = 32'h41C00000;
rContents[704] = 32'h18011005;
rContents[705] = 32'hD00FFEFE;
rContents[706] = 32'h183CC040;
rContents[707] = 32'h61C00000;
rContents[708] = 32'hD00FFED9;
rContents[709] = 32'h41C00000;
rContents[710] = 32'h61C00000;
rContents[711] = 32'h08CD0000;
rContents[712] = 32'h18DDCCFF;
rContents[713] = 32'h61D00000;
rContents[714] = 32'hD00FFED3;
rContents[715] = 32'h41D00000;
rContents[716] = 32'h18DDC8FF;
rContents[717] = 32'h61D00000;
rContents[718] = 32'hD00FFECF;
rContents[719] = 32'h41D00000;
rContents[720] = 32'h18DDC4FF;
rContents[721] = 32'h61D00000;
rContents[722] = 32'hD00FFECB;
rContents[723] = 32'h41D00000;
rContents[724] = 32'h18DDC0FF;
rContents[725] = 32'h61D00000;
rContents[726] = 32'hD00FFEC7;
rContents[727] = 32'h41D00000;
rContents[728] = 32'h41C00000;
rContents[729] = 32'h18E0C040;
rContents[730] = 32'h82000003;
rContents[731] = 32'h2D000095;
rContents[732] = 32'h80000006;
rContents[733] = 32'h18E0C048;
rContents[734] = 32'h82000003;
rContents[735] = 32'h2D000087;
rContents[736] = 32'h80000002;
rContents[737] = 32'h2D0000FF;
rContents[738] = 32'h61D00000;
rContents[739] = 32'hD00FFEBA;
rContents[740] = 32'h41D00000;
rContents[741] = 32'h2D00000A;
rContents[742] = 32'hD00FFED9;
rContents[743] = 32'h18E0F0FF;
rContents[744] = 32'h82000005;
rContents[745] = 32'h181DD001;
rContents[746] = 32'h18E0D000;
rContents[747] = 32'h81000002;
rContents[748] = 32'h800FFFFA;
rContents[749] = 32'h41D00000;
rContents[750] = 32'h41C00000;
rContents[751] = 32'hF0000000;
rContents[752] = 32'h61C00000;
rContents[753] = 32'h61D00000;
rContents[754] = 32'h61E00000;
rContents[755] = 32'h18111004;
rContents[756] = 32'h41D00000;
rContents[757] = 32'h41C00000;
rContents[758] = 32'h18011006;
rContents[759] = 32'h2F000001;
rContents[760] = 32'h61F00000;
rContents[761] = 32'hD00FFE90;
rContents[762] = 32'h41F00000;
rContents[763] = 32'h2F000011;
rContents[764] = 32'h61F00000;
rContents[765] = 32'h61D00000;
rContents[766] = 32'hD00FFFBD;
rContents[767] = 32'h18111002;
rContents[768] = 32'h18E0F000;
rContents[769] = 32'h8200001E;
rContents[770] = 32'hD00FFEBD;
rContents[771] = 32'h18E0F0FE;
rContents[772] = 32'h820FFFFE;
rContents[773] = 32'h2E000080;
rContents[774] = 32'h2D000000;
rContents[775] = 32'hD00FFEB8;
rContents[776] = 32'h186DF018;
rContents[777] = 32'hD00FFEB6;
rContents[778] = 32'h186FF010;
rContents[779] = 32'h103DDF00;
rContents[780] = 32'hD00FFEB3;
rContents[781] = 32'h186FF008;
rContents[782] = 32'h103DDF00;
rContents[783] = 32'hD00FFEB0;
rContents[784] = 32'h103DDF00;
rContents[785] = 32'h6CD00000;
rContents[786] = 32'h180CC001;
rContents[787] = 32'h181EE001;
rContents[788] = 32'h18E0E000;
rContents[789] = 32'h820FFFF2;
rContents[790] = 32'hD00FFEA9;
rContents[791] = 32'hD00FFEA8;
rContents[792] = 32'h2F000000;
rContents[793] = 32'h61F00000;
rContents[794] = 32'hD00FFE6F;
rContents[795] = 32'h41F00000;
rContents[796] = 32'hD00FFEA3;
rContents[797] = 32'h2F000000;
rContents[798] = 32'h80000006;
rContents[799] = 32'h2F000000;
rContents[800] = 32'h61F00000;
rContents[801] = 32'hD00FFE68;
rContents[802] = 32'h41F00000;
rContents[803] = 32'h2F0000FF;
rContents[804] = 32'h41E00000;
rContents[805] = 32'h41D00000;
rContents[806] = 32'h41C00000;
rContents[807] = 32'hF0000000;
rContents[808] = 32'h61C00000;
rContents[809] = 32'h61D00000;
rContents[810] = 32'h61E00000;
rContents[811] = 32'h18111004;
rContents[812] = 32'h41D00000;
rContents[813] = 32'h41C00000;
rContents[814] = 32'h18011006;
rContents[815] = 32'h2F000001;
rContents[816] = 32'h61F00000;
rContents[817] = 32'hD00FFE58;
rContents[818] = 32'h41F00000;
rContents[819] = 32'h2F000018;
rContents[820] = 32'h61F00000;
rContents[821] = 32'h61D00000;
rContents[822] = 32'hD00FFF85;
rContents[823] = 32'h18111002;
rContents[824] = 32'h18E0F000;
rContents[825] = 32'h8200002E;
rContents[826] = 32'h2F0000FE;
rContents[827] = 32'h61F00000;
rContents[828] = 32'hD00FFE61;
rContents[829] = 32'h41F00000;
rContents[830] = 32'h2E000080;
rContents[831] = 32'h4CD00000;
rContents[832] = 32'h61C00000;
rContents[833] = 32'h182CDCFF;
rContents[834] = 32'h188DD018;
rContents[835] = 32'h61D00000;
rContents[836] = 32'hD00FFE59;
rContents[837] = 32'h41D00000;
rContents[838] = 32'h182CD8FF;
rContents[839] = 32'h188DD010;
rContents[840] = 32'h61D00000;
rContents[841] = 32'hD00FFE54;
rContents[842] = 32'h41D00000;
rContents[843] = 32'h182CD4FF;
rContents[844] = 32'h188DD008;
rContents[845] = 32'h61D00000;
rContents[846] = 32'hD00FFE4F;
rContents[847] = 32'h41D00000;
rContents[848] = 32'h182CD0FF;
rContents[849] = 32'h61D00000;
rContents[850] = 32'hD00FFE4B;
rContents[851] = 32'h41D00000;
rContents[852] = 32'h41C00000;
rContents[853] = 32'h180CC001;
rContents[854] = 32'h181EE001;
rContents[855] = 32'h18E0E000;
rContents[856] = 32'h820FFFE7;
rContents[857] = 32'h2F0000FF;
rContents[858] = 32'h61F00000;
rContents[859] = 32'hD00FFE42;
rContents[860] = 32'hD00FFE41;
rContents[861] = 32'h41F00000;
rContents[862] = 32'hD00FFE61;
rContents[863] = 32'h18E0F0FF;
rContents[864] = 32'h820FFFFE;
rContents[865] = 32'h2F000000;
rContents[866] = 32'h61F00000;
rContents[867] = 32'hD00FFE26;
rContents[868] = 32'h41F00000;
rContents[869] = 32'h2F000000;
rContents[870] = 32'h80000006;
rContents[871] = 32'h2F000000;
rContents[872] = 32'h61F00000;
rContents[873] = 32'hD00FFE20;
rContents[874] = 32'h41F00000;
rContents[875] = 32'h2F0000FF;
rContents[876] = 32'h41E00000;
rContents[877] = 32'h41D00000;
rContents[878] = 32'h41C00000;
rContents[879] = 32'hF0000000;
rContents[880] = 32'h61C00000;
rContents[881] = 32'h61D00000;
rContents[882] = 32'h18111003;
rContents[883] = 32'h41C00000;
rContents[884] = 32'h18011004;
rContents[885] = 32'h2D001FE1;
rContents[886] = 32'h6DC00000;
rContents[887] = 32'h2D001FE0;
rContents[888] = 32'h2C000000;
rContents[889] = 32'h6DC00000;
rContents[890] = 32'h41D00000;
rContents[891] = 32'h41C00000;
rContents[892] = 32'hF0000000;
rContents[893] = 32'h61C00000;
rContents[894] = 32'h61D00000;
rContents[895] = 32'h2C000000;
rContents[896] = 32'h2D000000;
rContents[897] = 32'h2F001FE0;
rContents[898] = 32'h6FC00000;
rContents[899] = 32'h2F0000FF;
rContents[900] = 32'h61F00000;
rContents[901] = 32'h61D00000;
rContents[902] = 32'hD00FFD88;
rContents[903] = 32'h41D00000;
rContents[904] = 32'h41F00000;
rContents[905] = 32'h2F000080;
rContents[906] = 32'h100FFC00;
rContents[907] = 32'h61F00000;
rContents[908] = 32'h2F000000;
rContents[909] = 32'h61F00000;
rContents[910] = 32'hD00FFD80;
rContents[911] = 32'h41F00000;
rContents[912] = 32'h41F00000;
rContents[913] = 32'h180CC001;
rContents[914] = 32'h18E0C050;
rContents[915] = 32'h820FFFF6;
rContents[916] = 32'h2F0000FF;
rContents[917] = 32'h61F00000;
rContents[918] = 32'hD00FFD8F;
rContents[919] = 32'h08DF0000;
rContents[920] = 32'h41F00000;
rContents[921] = 32'h180DD050;
rContents[922] = 32'h18E0D2C8;
rContents[923] = 32'h81000008;
rContents[924] = 32'h2F0000FF;
rContents[925] = 32'h61F00000;
rContents[926] = 32'h61D00000;
rContents[927] = 32'hD00FFD6F;
rContents[928] = 32'h41D00000;
rContents[929] = 32'h41F00000;
rContents[930] = 32'h800FFFE7;
rContents[931] = 32'h2C000000;
rContents[932] = 32'h2D000000;
rContents[933] = 32'h2F0000FF;
rContents[934] = 32'h61F00000;
rContents[935] = 32'h61D00000;
rContents[936] = 32'hD00FFD66;
rContents[937] = 32'h41D00000;
rContents[938] = 32'h41F00000;
rContents[939] = 32'h41D00000;
rContents[940] = 32'h41C00000;
rContents[941] = 32'hF0000000;
rContents[942] = 32'h61C00000;
rContents[943] = 32'h61D00000;
rContents[944] = 32'h18111003;
rContents[945] = 32'h41D00000;
rContents[946] = 32'h41C00000;
rContents[947] = 32'h18011005;
rContents[948] = 32'h2F001FE0;
rContents[949] = 32'h6FC00000;
rContents[950] = 32'h186CD004;
rContents[951] = 32'h186DD006;
rContents[952] = 32'h100DDC00;
rContents[953] = 32'h2F0000FF;
rContents[954] = 32'h61F00000;
rContents[955] = 32'h61D00000;
rContents[956] = 32'hD00FFD52;
rContents[957] = 32'h41D00000;
rContents[958] = 32'h41F00000;
rContents[959] = 32'h41D00000;
rContents[960] = 32'h41C00000;
rContents[961] = 32'hF0000000;
rContents[962] = 32'hF0000000;
rContents[963] = 32'h61C00000;
rContents[964] = 32'h18111002;
rContents[965] = 32'h41C00000;
rContents[966] = 32'h18011003;
rContents[967] = 32'h18E0C020;
rContents[968] = 32'h8B00001B;
rContents[969] = 32'h18E0C00D;
rContents[970] = 32'h82000005;
rContents[971] = 32'h2C000000;
rContents[972] = 32'h2F001FE0;
rContents[973] = 32'h6FC00000;
rContents[974] = 32'h8000003A;
rContents[975] = 32'h18E0C00A;
rContents[976] = 32'h82000012;
rContents[977] = 32'h2F0000FF;
rContents[978] = 32'h61F00000;
rContents[979] = 32'hD00FFD52;
rContents[980] = 32'h08CF0000;
rContents[981] = 32'h41F00000;
rContents[982] = 32'h180CC050;
rContents[983] = 32'h18E0C2C8;
rContents[984] = 32'h82000003;
rContents[985] = 32'hD00FFFA4;
rContents[986] = 32'h8000002E;
rContents[987] = 32'h2F0000FF;
rContents[988] = 32'h61F00000;
rContents[989] = 32'h61C00000;
rContents[990] = 32'hD00FFD30;
rContents[991] = 32'h41C00000;
rContents[992] = 32'h41F00000;
rContents[993] = 32'h80000027;
rContents[994] = 32'h80000026;
rContents[995] = 32'h2F001FE0;
rContents[996] = 32'h4FF00000;
rContents[997] = 32'h180FF080;
rContents[998] = 32'h61F00000;
rContents[999] = 32'h2F001FE1;
rContents[1000] = 32'h4FF00000;
rContents[1001] = 32'h186FF008;
rContents[1002] = 32'h103CCF00;
rContents[1003] = 32'h61C00000;
rContents[1004] = 32'hD00FFD22;
rContents[1005] = 32'h41C00000;
rContents[1006] = 32'h41F00000;
rContents[1007] = 32'h2F001FE0;
rContents[1008] = 32'h4FC00000;
rContents[1009] = 32'h180CC001;
rContents[1010] = 32'h6FC00000;
rContents[1011] = 32'h18E0C050;
rContents[1012] = 32'h82000014;
rContents[1013] = 32'h2C000000;
rContents[1014] = 32'h2F001FE0;
rContents[1015] = 32'h6FC00000;
rContents[1016] = 32'h2F0000FF;
rContents[1017] = 32'h61F00000;
rContents[1018] = 32'hD00FFD2B;
rContents[1019] = 32'h08CF0000;
rContents[1020] = 32'h41F00000;
rContents[1021] = 32'h180CC050;
rContents[1022] = 32'h18E0C2C8;
rContents[1023] = 32'h81000008;
rContents[1024] = 32'h2F0000FF;
rContents[1025] = 32'h61F00000;
rContents[1026] = 32'h61C00000;
rContents[1027] = 32'hD00FFD0B;
rContents[1028] = 32'h41C00000;
rContents[1029] = 32'h41F00000;
rContents[1030] = 32'h80000002;
rContents[1031] = 32'hD00FFF76;
rContents[1032] = 32'h41C00000;
rContents[1033] = 32'hF0000000;
rContents[1034] = 32'h0A0A416E;
rContents[1035] = 32'h20657272;
rContents[1036] = 32'h6F722068;
rContents[1037] = 32'h6173206F;
rContents[1038] = 32'h63637572;
rContents[1039] = 32'h65642E0A;
rContents[1040] = 32'h00000000;
rContents[1041] = 32'h0A0A4120;
rContents[1042] = 32'h66617461;
rContents[1043] = 32'h6C206572;
rContents[1044] = 32'h726F7220;
rContents[1045] = 32'h68617320;
rContents[1046] = 32'h6F636375;
rContents[1047] = 32'h7265642E;
rContents[1048] = 32'h0A000000;
rContents[1049] = 32'h43616C6C;
rContents[1050] = 32'h65642061;
rContents[1051] = 32'h74200000;
rContents[1052] = 32'h53746163;
rContents[1053] = 32'h6B747261;
rContents[1054] = 32'h63652028;
rContents[1055] = 32'h746F7020;
rContents[1056] = 32'h3136293A;
rContents[1057] = 32'h0A000000;
rContents[1058] = 32'h52656769;
rContents[1059] = 32'h73746572;
rContents[1060] = 32'h733A0A00;
rContents[1061] = 32'h52657375;
rContents[1062] = 32'h6D696E67;
rContents[1063] = 32'h2E0A0A00;
rContents[1064] = 32'h48616C74;
rContents[1065] = 32'h696E672E;
rContents[1066] = 32'h0A0A0000;
rContents[1067] = 32'h80000001;
rContents[1068] = 32'h2F000411;
rContents[1069] = 32'h61F00000;
rContents[1070] = 32'hD00FFDDC;
rContents[1071] = 32'h41F00000;
rContents[1072] = 32'h2F000419;
rContents[1073] = 32'h61F00000;
rContents[1074] = 32'hD00FFDD8;
rContents[1075] = 32'h41F00000;
rContents[1076] = 32'hD00FFDA9;
rContents[1077] = 32'h04200000;
rContents[1078] = 32'h61F00000;
rContents[1079] = 32'h2F000419;
rContents[1080] = 32'h61F00000;
rContents[1081] = 32'hD00FFDD1;
rContents[1082] = 32'h41F00000;
rContents[1083] = 32'h2F0000F0;
rContents[1084] = 32'h181FF001;
rContents[1085] = 32'h18E0F000;
rContents[1086] = 32'h820FFFFE;
rContents[1087] = 32'h18111001;
rContents[1088] = 32'hD00FFD9D;
rContents[1089] = 32'h18011001;
rContents[1090] = 32'h2F00000A;
rContents[1091] = 32'h61F00000;
rContents[1092] = 32'hD0000013;
rContents[1093] = 32'h41F00000;
rContents[1094] = 32'h2F00000D;
rContents[1095] = 32'h61F00000;
rContents[1096] = 32'hD000000F;
rContents[1097] = 32'h41F00000;
rContents[1098] = 32'h41F00000;
rContents[1099] = 32'hF0000000;
rContents[1100] = 32'hF0000000;
rContents[1101] = 32'hF0000000;
rContents[1102] = 32'h4C656D6F;
rContents[1103] = 32'h6E207630;
rContents[1104] = 32'h2E32202D;
rContents[1105] = 32'h20666F72;
rContents[1106] = 32'h20657052;
rContents[1107] = 32'h49534320;
rContents[1108] = 32'h76352073;
rContents[1109] = 32'h79737465;
rContents[1110] = 32'h6D730000;
rContents[1111] = 32'h800FFCEA;
rContents[1112] = 32'h800FFD05;
rContents[1113] = 32'h800FFD84;
rContents[1114] = 32'h800FFDB0;
rContents[1115] = 32'h800FFFD1;
rContents[1116] = 32'h210017FF;
rContents[1117] = 32'h2800044E;
rContents[1118] = 32'h61800000;
rContents[1119] = 32'hD00FFFFB;
rContents[1120] = 32'h41800000;
rContents[1121] = 32'h26001000;
rContents[1122] = 32'h29000000;
rContents[1123] = 32'h2800000A;
rContents[1124] = 32'h61800000;
rContents[1125] = 32'hD00FFFF2;
rContents[1126] = 32'h41800000;
rContents[1127] = 32'h2800000D;
rContents[1128] = 32'h61800000;
rContents[1129] = 32'hD00FFFEE;
rContents[1130] = 32'h41800000;
rContents[1131] = 32'h2800003E;
rContents[1132] = 32'h61800000;
rContents[1133] = 32'hD00FFFEA;
rContents[1134] = 32'h41800000;
rContents[1135] = 32'hD00FFFE9;
rContents[1136] = 32'h18E0F008;
rContents[1137] = 32'h8200000E;
rContents[1138] = 32'h18E06000;
rContents[1139] = 32'h82000002;
rContents[1140] = 32'h800FFFFB;
rContents[1141] = 32'h18166002;
rContents[1142] = 32'h18199001;
rContents[1143] = 32'h46F00000;
rContents[1144] = 32'h61F00000;
rContents[1145] = 32'hD00FFFDE;
rContents[1146] = 32'h41F00000;
rContents[1147] = 32'h18066001;
rContents[1148] = 32'h2F000000;
rContents[1149] = 32'h66F00000;
rContents[1150] = 32'h800FFFF1;
rContents[1151] = 32'h18E0F00D;
rContents[1152] = 32'h82000003;
rContents[1153] = 32'h66F00000;
rContents[1154] = 32'h8000000A;
rContents[1155] = 32'h18F09180;
rContents[1156] = 32'h820FFFEB;
rContents[1157] = 32'h61F00000;
rContents[1158] = 32'hD00FFFD1;
rContents[1159] = 32'h41F00000;
rContents[1160] = 32'h66F00000;
rContents[1161] = 32'h18066001;
rContents[1162] = 32'h18099001;
rContents[1163] = 32'h800FFFE4;
rContents[1164] = 32'h26001000;
rContents[1165] = 32'h27000000;
rContents[1166] = 32'h46900000;
rContents[1167] = 32'h18E0900D;
rContents[1168] = 32'h82000005;
rContents[1169] = 32'h18E0703A;
rContents[1170] = 32'h82000002;
rContents[1171] = 32'h41800000;
rContents[1172] = 32'h800FFFCD;
rContents[1173] = 32'h18E09052;
rContents[1174] = 32'h8200000C;
rContents[1175] = 32'h2800000A;
rContents[1176] = 32'h61800000;
rContents[1177] = 32'hD00FFFBE;
rContents[1178] = 32'h41800000;
rContents[1179] = 32'h2800000D;
rContents[1180] = 32'h61800000;
rContents[1181] = 32'hD00FFFBA;
rContents[1182] = 32'h41800000;
rContents[1183] = 32'hD0400000;
rContents[1184] = 32'h18066001;
rContents[1185] = 32'h800FFFED;
rContents[1186] = 32'h18E0903A;
rContents[1187] = 32'h82000005;
rContents[1188] = 32'h2700003A;
rContents[1189] = 32'h61400000;
rContents[1190] = 32'h18066001;
rContents[1191] = 32'h800FFFE7;
rContents[1192] = 32'h18E0902E;
rContents[1193] = 32'h82000007;
rContents[1194] = 32'h18E0703A;
rContents[1195] = 32'h82000002;
rContents[1196] = 32'h41800000;
rContents[1197] = 32'h2700002E;
rContents[1198] = 32'h18066001;
rContents[1199] = 32'h800FFFDF;
rContents[1200] = 32'h18E09020;
rContents[1201] = 32'h82000003;
rContents[1202] = 32'h18066001;
rContents[1203] = 32'h800FFFDB;
rContents[1204] = 32'h25000000;
rContents[1205] = 32'h46900000;
rContents[1206] = 32'h18199030;
rContents[1207] = 32'h18E0900A;
rContents[1208] = 32'h84000007;
rContents[1209] = 32'h18199007;
rContents[1210] = 32'h18E0900A;
rContents[1211] = 32'h84000008;
rContents[1212] = 32'h18E09010;
rContents[1213] = 32'h84000002;
rContents[1214] = 32'h80000005;
rContents[1215] = 32'h18655004;
rContents[1216] = 32'h10355900;
rContents[1217] = 32'h18066001;
rContents[1218] = 32'h800FFFF3;
rContents[1219] = 32'h46900000;
rContents[1220] = 32'h18E0703A;
rContents[1221] = 32'h82000004;
rContents[1222] = 32'h64500000;
rContents[1223] = 32'h18044001;
rContents[1224] = 32'h800FFFC6;
rContents[1225] = 32'h61400000;
rContents[1226] = 32'h08450000;
rContents[1227] = 32'h18E0902E;
rContents[1228] = 32'h82000003;
rContents[1229] = 32'h41800000;
rContents[1230] = 32'h800FFFC0;
rContents[1231] = 32'h18E07000;
rContents[1232] = 32'h8200001A;
rContents[1233] = 32'h41800000;
rContents[1234] = 32'h2800000A;
rContents[1235] = 32'h61800000;
rContents[1236] = 32'hD00FFF83;
rContents[1237] = 32'h41800000;
rContents[1238] = 32'h2800000D;
rContents[1239] = 32'h61800000;
rContents[1240] = 32'hD00FFF7F;
rContents[1241] = 32'h41800000;
rContents[1242] = 32'h61400000;
rContents[1243] = 32'hD00FFD02;
rContents[1244] = 32'h41400000;
rContents[1245] = 32'h2800003A;
rContents[1246] = 32'h61800000;
rContents[1247] = 32'hD00FFF78;
rContents[1248] = 32'h41800000;
rContents[1249] = 32'h28000020;
rContents[1250] = 32'h61800000;
rContents[1251] = 32'hD00FFF74;
rContents[1252] = 32'h41800000;
rContents[1253] = 32'h44800000;
rContents[1254] = 32'h61800000;
rContents[1255] = 32'hD00FFF72;
rContents[1256] = 32'h41800000;
rContents[1257] = 32'h800FFFA5;
rContents[1258] = 32'h18E0702E;
rContents[1259] = 32'hD20FFF70;
rContents[1260] = 32'h08840000;
rContents[1261] = 32'h41400000;
rContents[1262] = 32'h10E08400;
rContents[1263] = 32'h8B000002;
rContents[1264] = 32'h08840000;
rContents[1265] = 32'h101A8400;
rContents[1266] = 32'h180AA001;
rContents[1267] = 32'h61400000;
rContents[1268] = 32'h2800000A;
rContents[1269] = 32'h61800000;
rContents[1270] = 32'hD00FFF61;
rContents[1271] = 32'h41800000;
rContents[1272] = 32'h2800000D;
rContents[1273] = 32'h61800000;
rContents[1274] = 32'hD00FFF5D;
rContents[1275] = 32'h41800000;
rContents[1276] = 32'h61400000;
rContents[1277] = 32'hD00FFCE0;
rContents[1278] = 32'h41400000;
rContents[1279] = 32'h2800003A;
rContents[1280] = 32'h61800000;
rContents[1281] = 32'hD00FFF56;
rContents[1282] = 32'h41800000;
rContents[1283] = 32'h18E0A008;
rContents[1284] = 32'h83000003;
rContents[1285] = 32'h08BA0000;
rContents[1286] = 32'h80000002;
rContents[1287] = 32'h2B000008;
rContents[1288] = 32'h101AAB00;
rContents[1289] = 32'h28000020;
rContents[1290] = 32'h61800000;
rContents[1291] = 32'hD00FFF4C;
rContents[1292] = 32'h41800000;
rContents[1293] = 32'h44800000;
rContents[1294] = 32'h61800000;
rContents[1295] = 32'hD00FFF4A;
rContents[1296] = 32'h41800000;
rContents[1297] = 32'h18044001;
rContents[1298] = 32'h181BB001;
rContents[1299] = 32'h18E0B000;
rContents[1300] = 32'h820FFFF5;
rContents[1301] = 32'h18E0A000;
rContents[1302] = 32'h820FFFDE;
rContents[1303] = 32'h41400000;
rContents[1304] = 32'h27000000;
rContents[1305] = 32'h800FFF75;
    end

endmodule

/*  Program 1 - square wave generator over GPIO
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808000;
        rContents[8] = 32'h3500FFFF;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25000000;
        rContents[17] = 32'h08650000;
        rContents[18] = 32'h36808002;
        rContents[19] = 32'h64600001;
        rContents[20] = 32'h27010005;
        rContents[21] = 32'h64700000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h04000000;
        rContents[26] = 32'h18B5580F;
        rContents[27] = 32'h18055001;
        rContents[28] = 32'h800FFFF5;
        rContents[29] = 32'h0;
        rContents[30] = 32'h0;
        rContents[31] = 32'h0;
        rContents[32] = 32'h0;
        rContents[33] = 32'h0;
        rContents[34] = 32'h0;
        rContents[35] = 32'h0; */
        
/*  Program 2 - print some 'H's over the serial link
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808101;
        rContents[8] = 32'h35000048;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25808100;
        rContents[17] = 32'h35000080;
        rContents[18] = 32'h64500001;
        rContents[19] = 32'h27010005;
        rContents[20] = 32'h64700000;
        rContents[21] = 32'h04000000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h800FFFED; */
