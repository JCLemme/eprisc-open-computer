module epRISC_embeddedROM(iClk, iAddr, oData, iEnable);

    input iClk, iEnable;
    input [11:0] iAddr;
    output wire [31:0] oData;
    
    reg [31:0] rDataOut, rContents[0:4095];
    
    assign oData = (iEnable) ? rDataOut : 32'bz;
    
    always @(posedge iClk) begin
        rDataOut = rContents[iAddr];
    end
    
    initial begin
rContents[0] = 32'h8000001F;
rContents[1] = 32'h43F01FF0;
rContents[2] = 32'h61F00000;
rContents[3] = 32'hD000026E;
rContents[4] = 32'h63F01FF1;
rContents[5] = 32'h41F00000;
rContents[6] = 32'hF0000000;
rContents[7] = 32'hD000028C;
rContents[8] = 32'h63F01FF1;
rContents[9] = 32'hF0000000;
rContents[10] = 32'h43F01FF2;
rContents[11] = 32'h61F00000;
rContents[12] = 32'h43F01FF3;
rContents[13] = 32'h61F00000;
rContents[14] = 32'hD00003BD;
rContents[15] = 32'h63F01FF4;
rContents[16] = 32'h41F00000;
rContents[17] = 32'h41F00000;
rContents[18] = 32'hF0000000;
rContents[19] = 32'h43F01FF2;
rContents[20] = 32'h61F00000;
rContents[21] = 32'h43F01FF3;
rContents[22] = 32'h61F00000;
rContents[23] = 32'hD00003E9;
rContents[24] = 32'h63F01FF4;
rContents[25] = 32'h41F00000;
rContents[26] = 32'h41F00000;
rContents[27] = 32'hF0000000;
rContents[28] = 32'hD0000314;
rContents[29] = 32'h63F01FF5;
rContents[30] = 32'hF0000000;
rContents[31] = 32'h21001100;
rContents[32] = 32'h23000000;
rContents[33] = 32'hD00001B4;
rContents[34] = 32'h24007FFF;
rContents[35] = 32'h61400000;
rContents[36] = 32'h24000000;
rContents[37] = 32'h61400000;
rContents[38] = 32'hD00001BC;
rContents[39] = 32'h41400000;
rContents[40] = 32'h41400000;
rContents[41] = 32'hD0000460;
rContents[42] = 32'h24000117;
rContents[43] = 32'h61400000;
rContents[44] = 32'hD00002D3;
rContents[45] = 32'h41400000;
rContents[46] = 32'h2400019E;
rContents[47] = 32'h61400000;
rContents[48] = 32'hD00002CF;
rContents[49] = 32'h41400000;
rContents[50] = 32'h240001C0;
rContents[51] = 32'h61400000;
rContents[52] = 32'hD00002CB;
rContents[53] = 32'h41400000;
rContents[54] = 32'h24000041;
rContents[55] = 32'h61400000;
rContents[56] = 32'hD0000239;
rContents[57] = 32'h41400000;
rContents[58] = 32'h24000128;
rContents[59] = 32'h61400000;
rContents[60] = 32'hD00002C3;
rContents[61] = 32'h41400000;
rContents[62] = 32'hD00002F2;
rContents[63] = 32'h61F00000;
rContents[64] = 32'h24000147;
rContents[65] = 32'h18E0F0FF;
rContents[66] = 32'h81000002;
rContents[67] = 32'h2400013E;
rContents[68] = 32'h61400000;
rContents[69] = 32'hD00002BA;
rContents[70] = 32'h41400000;
rContents[71] = 32'h41F00000;
rContents[72] = 32'h18E0F0FF;
rContents[73] = 32'h810000C9;
rContents[74] = 32'h2400014F;
rContents[75] = 32'h61400000;
rContents[76] = 32'hD00002B3;
rContents[77] = 32'h41400000;
rContents[78] = 32'h24003000;
rContents[79] = 32'h61400000;
rContents[80] = 32'h24000000;
rContents[81] = 32'h61400000;
rContents[82] = 32'hD00003AE;
rContents[83] = 32'h41400000;
rContents[84] = 32'h41400000;
rContents[85] = 32'h24003000;
rContents[86] = 32'h44F00000;
rContents[87] = 32'h18E0FCEA;
rContents[88] = 32'h81000006;
rContents[89] = 32'h24000155;
rContents[90] = 32'h61400000;
rContents[91] = 32'hD00002A4;
rContents[92] = 32'h41400000;
rContents[93] = 32'h800000B5;
rContents[94] = 32'h2400015E;
rContents[95] = 32'h61400000;
rContents[96] = 32'hD000029F;
rContents[97] = 32'h41400000;
rContents[98] = 32'h24003001;
rContents[99] = 32'h61400000;
rContents[100] = 32'h2400000C;
rContents[101] = 32'h61400000;
rContents[102] = 32'hD00002AF;
rContents[103] = 32'h41400000;
rContents[104] = 32'h41400000;
rContents[105] = 32'h24000162;
rContents[106] = 32'h61400000;
rContents[107] = 32'hD0000294;
rContents[108] = 32'h41400000;
rContents[109] = 32'h24003000;
rContents[110] = 32'h44F00000;
rContents[111] = 32'h18E0F000;
rContents[112] = 32'h82000006;
rContents[113] = 32'h24000166;
rContents[114] = 32'h61400000;
rContents[115] = 32'hD000028C;
rContents[116] = 32'h41400000;
rContents[117] = 32'h8000009D;
rContents[118] = 32'h2400016E;
rContents[119] = 32'h61400000;
rContents[120] = 32'hD0000287;
rContents[121] = 32'h41400000;
rContents[122] = 32'h24003004;
rContents[123] = 32'h44F00000;
rContents[124] = 32'h61F00000;
rContents[125] = 32'h24000002;
rContents[126] = 32'h61400000;
rContents[127] = 32'hD000024B;
rContents[128] = 32'h41400000;
rContents[129] = 32'h41F00000;
rContents[130] = 32'h24000171;
rContents[131] = 32'h61400000;
rContents[132] = 32'hD000027B;
rContents[133] = 32'h41400000;
rContents[134] = 32'h24000177;
rContents[135] = 32'h61400000;
rContents[136] = 32'hD0000277;
rContents[137] = 32'h41400000;
rContents[138] = 32'h24003004;
rContents[139] = 32'h44600000;
rContents[140] = 32'h18656002;
rContents[141] = 32'h18666001;
rContents[142] = 32'h10066500;
rContents[143] = 32'h25003005;
rContents[144] = 32'h10065600;
rContents[145] = 32'h27000000;
rContents[146] = 32'h240001D4;
rContents[147] = 32'h61400000;
rContents[148] = 32'hD000026B;
rContents[149] = 32'h41400000;
rContents[150] = 32'h61700000;
rContents[151] = 32'h24000002;
rContents[152] = 32'h61400000;
rContents[153] = 32'hD0000231;
rContents[154] = 32'h41400000;
rContents[155] = 32'h41700000;
rContents[156] = 32'h2400017D;
rContents[157] = 32'h61400000;
rContents[158] = 32'hD0000261;
rContents[159] = 32'h41400000;
rContents[160] = 32'h61500000;
rContents[161] = 32'h2400000C;
rContents[162] = 32'h61400000;
rContents[163] = 32'hD0000272;
rContents[164] = 32'h41400000;
rContents[165] = 32'h41500000;
rContents[166] = 32'h18055003;
rContents[167] = 32'h24000180;
rContents[168] = 32'h61400000;
rContents[169] = 32'hD0000256;
rContents[170] = 32'h41400000;
rContents[171] = 32'h45400000;
rContents[172] = 32'h61400000;
rContents[173] = 32'hD0000204;
rContents[174] = 32'h41400000;
rContents[175] = 32'h18055001;
rContents[176] = 32'h24000183;
rContents[177] = 32'h61400000;
rContents[178] = 32'hD000024D;
rContents[179] = 32'h41400000;
rContents[180] = 32'h45400000;
rContents[181] = 32'h61400000;
rContents[182] = 32'hD00001FB;
rContents[183] = 32'h41400000;
rContents[184] = 32'h18055001;
rContents[185] = 32'h24000186;
rContents[186] = 32'h61400000;
rContents[187] = 32'hD0000244;
rContents[188] = 32'h41400000;
rContents[189] = 32'h45400000;
rContents[190] = 32'h61400000;
rContents[191] = 32'hD00001F2;
rContents[192] = 32'h41400000;
rContents[193] = 32'h18055001;
rContents[194] = 32'h240001D3;
rContents[195] = 32'h61400000;
rContents[196] = 32'hD000023B;
rContents[197] = 32'h41400000;
rContents[198] = 32'h18077001;
rContents[199] = 32'h10E05600;
rContents[200] = 32'h840FFFCA;
rContents[201] = 32'h240001D3;
rContents[202] = 32'h61400000;
rContents[203] = 32'hD0000234;
rContents[204] = 32'h41400000;
rContents[205] = 32'h24000188;
rContents[206] = 32'h61400000;
rContents[207] = 32'hD0000230;
rContents[208] = 32'h41400000;
rContents[209] = 32'hD0000160;
rContents[210] = 32'h61F00000;
rContents[211] = 32'hD0000142;
rContents[212] = 32'hD0000412;
rContents[213] = 32'h41F00000;
rContents[214] = 32'h18E0F047;
rContents[215] = 32'h8300000E;
rContents[216] = 32'h181FF030;
rContents[217] = 32'h18E0F00A;
rContents[218] = 32'h84000014;
rContents[219] = 32'h181FF007;
rContents[220] = 32'h18E0F00A;
rContents[221] = 32'h84000003;
rContents[222] = 32'h18E0F010;
rContents[223] = 32'h8400000F;
rContents[224] = 32'h240001D3;
rContents[225] = 32'h61400000;
rContents[226] = 32'hD000021D;
rContents[227] = 32'h41400000;
rContents[228] = 32'h800FFFE9;
rContents[229] = 32'h61F00000;
rContents[230] = 32'h240001D3;
rContents[231] = 32'h61400000;
rContents[232] = 32'hD0000217;
rContents[233] = 32'h41400000;
rContents[234] = 32'h41F00000;
rContents[235] = 32'h18E0F04D;
rContents[236] = 32'h81000026;
rContents[237] = 32'h800FFFE0;
rContents[238] = 32'h240001D3;
rContents[239] = 32'h61400000;
rContents[240] = 32'hD000020F;
rContents[241] = 32'h41400000;
rContents[242] = 32'h61F00000;
rContents[243] = 32'h24000198;
rContents[244] = 32'h61400000;
rContents[245] = 32'hD000020A;
rContents[246] = 32'h41400000;
rContents[247] = 32'h41F00000;
rContents[248] = 32'h1865F002;
rContents[249] = 32'h186FF001;
rContents[250] = 32'h100FF500;
rContents[251] = 32'h25003005;
rContents[252] = 32'h10085F00;
rContents[253] = 32'h48500003;
rContents[254] = 32'h48600004;
rContents[255] = 32'h48700005;
rContents[256] = 32'h61700000;
rContents[257] = 32'h61500000;
rContents[258] = 32'hD00002FE;
rContents[259] = 32'h41500000;
rContents[260] = 32'h41700000;
rContents[261] = 32'h18E0F000;
rContents[262] = 32'h8200000C;
rContents[263] = 32'h18055001;
rContents[264] = 32'h18077080;
rContents[265] = 32'h18166001;
rContents[266] = 32'h18E06000;
rContents[267] = 32'h820FFFF5;
rContents[268] = 32'hD0000396;
rContents[269] = 32'h48700005;
rContents[270] = 32'h61700000;
rContents[271] = 32'hD00001A2;
rContents[272] = 32'h41700000;
rContents[273] = 32'h80700000;
rContents[274] = 32'h240001CD;
rContents[275] = 32'h61400000;
rContents[276] = 32'hD00001EB;
rContents[277] = 32'h41400000;
rContents[278] = 32'h80000486;
rContents[279] = 32'h65705249;
rContents[280] = 32'h53432042;
rContents[281] = 32'h6F6F746C;
rContents[282] = 32'h6F616465;
rContents[283] = 32'h72207633;
rContents[284] = 32'h2E340A0D;
rContents[285] = 32'h636F7079;
rContents[286] = 32'h72696768;
rContents[287] = 32'h74203230;
rContents[288] = 32'h31352D32;
rContents[289] = 32'h30313720;
rContents[290] = 32'h50726F70;
rContents[291] = 32'h6F727469;
rContents[292] = 32'h6F6E616C;
rContents[293] = 32'h204C6162;
rContents[294] = 32'h730A0D0A;
rContents[295] = 32'h0D000000;
rContents[296] = 32'h41747465;
rContents[297] = 32'h6D707469;
rContents[298] = 32'h6E672074;
rContents[299] = 32'h6F206D6F;
rContents[300] = 32'h756E7420;
rContents[301] = 32'h53442063;
rContents[302] = 32'h61726420;
rContents[303] = 32'h696E2073;
rContents[304] = 32'h6C6F7420;
rContents[305] = 32'h412E2E2E;
rContents[306] = 32'h0A0D0000;
rContents[307] = 32'h41747465;
rContents[308] = 32'h6D707469;
rContents[309] = 32'h6E672074;
rContents[310] = 32'h6F206D6F;
rContents[311] = 32'h756E7420;
rContents[312] = 32'h53442063;
rContents[313] = 32'h61726420;
rContents[314] = 32'h696E2073;
rContents[315] = 32'h6C6F7420;
rContents[316] = 32'h422E2E2E;
rContents[317] = 32'h0A0D0000;
rContents[318] = 32'h20205344;
rContents[319] = 32'h20636172;
rContents[320] = 32'h64206D6F;
rContents[321] = 32'h756E7465;
rContents[322] = 32'h64207375;
rContents[323] = 32'h63636573;
rContents[324] = 32'h7366756C;
rContents[325] = 32'h6C792E0A;
rContents[326] = 32'h0D0A0D00;
rContents[327] = 32'h20204572;
rContents[328] = 32'h726F7220;
rContents[329] = 32'h6D6F756E;
rContents[330] = 32'h74696E67;
rContents[331] = 32'h20534420;
rContents[332] = 32'h63617264;
rContents[333] = 32'h2E0A0D0A;
rContents[334] = 32'h0D000000;
rContents[335] = 32'h46657463;
rContents[336] = 32'h68696E67;
rContents[337] = 32'h20646973;
rContents[338] = 32'h6B20696E;
rContents[339] = 32'h666F2E2E;
rContents[340] = 32'h2E0A0D00;
rContents[341] = 32'h20204469;
rContents[342] = 32'h736B2061;
rContents[343] = 32'h70706561;
rContents[344] = 32'h72732074;
rContents[345] = 32'h6F206265;
rContents[346] = 32'h20636F72;
rContents[347] = 32'h72757074;
rContents[348] = 32'h2E0A0D0A;
rContents[349] = 32'h0D000000;
rContents[350] = 32'h2020466F;
rContents[351] = 32'h756E6420;
rContents[352] = 32'h6469736B;
rContents[353] = 32'h20270000;
rContents[354] = 32'h27206174;
rContents[355] = 32'h20626C6F;
rContents[356] = 32'h636B2030;
rContents[357] = 32'h2E0A0D00;
rContents[358] = 32'h20204469;
rContents[359] = 32'h736B2061;
rContents[360] = 32'h70706561;
rContents[361] = 32'h72732074;
rContents[362] = 32'h6F206265;
rContents[363] = 32'h20656D70;
rContents[364] = 32'h74792E0A;
rContents[365] = 32'h0D0A0D00;
rContents[366] = 32'h2020466F;
rContents[367] = 32'h756E6420;
rContents[368] = 32'h00000000;
rContents[369] = 32'h20656E74;
rContents[370] = 32'h72696573;
rContents[371] = 32'h206F6E20;
rContents[372] = 32'h6469736B;
rContents[373] = 32'h2E0A0D0A;
rContents[374] = 32'h0D000000;
rContents[375] = 32'h41766169;
rContents[376] = 32'h6C61626C;
rContents[377] = 32'h6520656E;
rContents[378] = 32'h74726965;
rContents[379] = 32'h733A0A0D;
rContents[380] = 32'h00000000;
rContents[381] = 32'h3A20456E;
rContents[382] = 32'h74727920;
rContents[383] = 32'h27000000;
rContents[384] = 32'h273A2073;
rContents[385] = 32'h74617274;
rContents[386] = 32'h20000000;
rContents[387] = 32'h2C206C65;
rContents[388] = 32'h6E677468;
rContents[389] = 32'h20000000;
rContents[390] = 32'h2C206C6F;
rContents[391] = 32'h61642000;
rContents[392] = 32'h53656C65;
rContents[393] = 32'h63742061;
rContents[394] = 32'h6E20656E;
rContents[395] = 32'h74727920;
rContents[396] = 32'h746F2065;
rContents[397] = 32'h78656375;
rContents[398] = 32'h74652C20;
rContents[399] = 32'h6F722074;
rContents[400] = 32'h79706520;
rContents[401] = 32'h274D2720;
rContents[402] = 32'h746F2065;
rContents[403] = 32'h6E746572;
rContents[404] = 32'h20746865;
rContents[405] = 32'h206D6F6E;
rContents[406] = 32'h69746F72;
rContents[407] = 32'h3A200000;
rContents[408] = 32'h20204C6F;
rContents[409] = 32'h6164696E;
rContents[410] = 32'h6720656E;
rContents[411] = 32'h7472792E;
rContents[412] = 32'h2E2E0A0D;
rContents[413] = 32'h0A0D0000;
rContents[414] = 32'h53746172;
rContents[415] = 32'h74696E67;
rContents[416] = 32'h20504F53;
rContents[417] = 32'h54732E2E;
rContents[418] = 32'h2E0A0D00;
rContents[419] = 32'h20204D65;
rContents[420] = 32'h6D6F7279;
rContents[421] = 32'h20202020;
rContents[422] = 32'h20202020;
rContents[423] = 32'h20200000;
rContents[424] = 32'h20205541;
rContents[425] = 32'h52542020;
rContents[426] = 32'h20202020;
rContents[427] = 32'h20202020;
rContents[428] = 32'h20200000;
rContents[429] = 32'h20205350;
rContents[430] = 32'h49202020;
rContents[431] = 32'h20202020;
rContents[432] = 32'h20202020;
rContents[433] = 32'h20200000;
rContents[434] = 32'h20207379;
rContents[435] = 32'h73582042;
rContents[436] = 32'h75732020;
rContents[437] = 32'h20202020;
rContents[438] = 32'h20200000;
rContents[439] = 32'h2020492F;
rContents[440] = 32'h4F20436F;
rContents[441] = 32'h6E74726F;
rContents[442] = 32'h6C6C6572;
rContents[443] = 32'h20200000;
rContents[444] = 32'h4F4B0A0D;
rContents[445] = 32'h00000000;
rContents[446] = 32'h4641494C;
rContents[447] = 32'h0A0D0000;
rContents[448] = 32'h2020504F;
rContents[449] = 32'h53542073;
rContents[450] = 32'h75636365;
rContents[451] = 32'h73736675;
rContents[452] = 32'h6C2E0A0D;
rContents[453] = 32'h0A0D0000;
rContents[454] = 32'h2020504F;
rContents[455] = 32'h53542075;
rContents[456] = 32'h6E737563;
rContents[457] = 32'h63657373;
rContents[458] = 32'h66756C2E;
rContents[459] = 32'h0A0D0A0D;
rContents[460] = 32'h00000000;
rContents[461] = 32'h456E7465;
rContents[462] = 32'h72696E67;
rContents[463] = 32'h206D6F6E;
rContents[464] = 32'h69746F72;
rContents[465] = 32'h2E2E2E0A;
rContents[466] = 32'h0D0A0D00;
rContents[467] = 32'h0A0D0000;
rContents[468] = 32'h20200000;
rContents[469] = 32'h61C00000;
rContents[470] = 32'h2C002000;
rContents[471] = 32'h2F010001;
rContents[472] = 32'h6CF00000;
rContents[473] = 32'h04000000;
rContents[474] = 32'h04000000;
rContents[475] = 32'h04000000;
rContents[476] = 32'h04000000;
rContents[477] = 32'h4CF00000;
rContents[478] = 32'h18F0F001;
rContents[479] = 32'h820FFFFE;
rContents[480] = 32'h41C00000;
rContents[481] = 32'hF0000000;
rContents[482] = 32'h61E00000;
rContents[483] = 32'h61D00000;
rContents[484] = 32'h61C00000;
rContents[485] = 32'h18111004;
rContents[486] = 32'h2C002000;
rContents[487] = 32'h41D00000;
rContents[488] = 32'h41E00000;
rContents[489] = 32'h18011006;
rContents[490] = 32'h2F600008;
rContents[491] = 32'h103FFE00;
rContents[492] = 32'h186FF010;
rContents[493] = 32'h103FFD00;
rContents[494] = 32'h6CF00001;
rContents[495] = 32'h2F010005;
rContents[496] = 32'h6CF00000;
rContents[497] = 32'h4CF00000;
rContents[498] = 32'h18F0F001;
rContents[499] = 32'h820FFFFE;
rContents[500] = 32'h4CF00002;
rContents[501] = 32'h41C00000;
rContents[502] = 32'h41D00000;
rContents[503] = 32'h41E00000;
rContents[504] = 32'hF0000000;
rContents[505] = 32'h61E00000;
rContents[506] = 32'h61C00000;
rContents[507] = 32'h18111003;
rContents[508] = 32'h2C002000;
rContents[509] = 32'h41E00000;
rContents[510] = 32'h18011004;
rContents[511] = 32'h2F600000;
rContents[512] = 32'h103FFE00;
rContents[513] = 32'h186FF010;
rContents[514] = 32'h6CF00001;
rContents[515] = 32'h2F010005;
rContents[516] = 32'h6CF00000;
rContents[517] = 32'h4CF00000;
rContents[518] = 32'h18F0F001;
rContents[519] = 32'h820FFFFE;
rContents[520] = 32'h2F600000;
rContents[521] = 32'h103FFE00;
rContents[522] = 32'h186FF010;
rContents[523] = 32'h6CF00001;
rContents[524] = 32'h2F010005;
rContents[525] = 32'h6CF00000;
rContents[526] = 32'h4CF00000;
rContents[527] = 32'h18F0F001;
rContents[528] = 32'h820FFFFE;
rContents[529] = 32'h4CF00002;
rContents[530] = 32'h41C00000;
rContents[531] = 32'h41E00000;
rContents[532] = 32'hF0000000;
rContents[533] = 32'h61D00000;
rContents[534] = 32'h61C00000;
rContents[535] = 32'h18111003;
rContents[536] = 32'h2C002000;
rContents[537] = 32'h41D00000;
rContents[538] = 32'h18011004;
rContents[539] = 32'h2F000011;
rContents[540] = 32'h61F00000;
rContents[541] = 32'h61D00000;
rContents[542] = 32'hD00FFFC4;
rContents[543] = 32'h41D00000;
rContents[544] = 32'h41F00000;
rContents[545] = 32'h2F000010;
rContents[546] = 32'h61F00000;
rContents[547] = 32'h2F000080;
rContents[548] = 32'h61F00000;
rContents[549] = 32'hD00FFFBD;
rContents[550] = 32'h41D00000;
rContents[551] = 32'h41F00000;
rContents[552] = 32'h2F000010;
rContents[553] = 32'h61F00000;
rContents[554] = 32'hD00FFFCF;
rContents[555] = 32'h18F0F080;
rContents[556] = 32'h820FFFFE;
rContents[557] = 32'h41F00000;
rContents[558] = 32'h41C00000;
rContents[559] = 32'h41D00000;
rContents[560] = 32'hF0000000;
rContents[561] = 32'h61C00000;
rContents[562] = 32'h2C002000;
rContents[563] = 32'h2F808010;
rContents[564] = 32'h3F000020;
rContents[565] = 32'h6CF00001;
rContents[566] = 32'h2F010005;
rContents[567] = 32'h6CF00000;
rContents[568] = 32'h4CF00000;
rContents[569] = 32'h18F0F001;
rContents[570] = 32'h820FFFFE;
rContents[571] = 32'h2F800010;
rContents[572] = 32'h6CF00001;
rContents[573] = 32'h2F010005;
rContents[574] = 32'h6CF00000;
rContents[575] = 32'h4CF00000;
rContents[576] = 32'h18F0F001;
rContents[577] = 32'h820FFFFE;
rContents[578] = 32'h2F800010;
rContents[579] = 32'h6CF00001;
rContents[580] = 32'h2F010005;
rContents[581] = 32'h6CF00000;
rContents[582] = 32'h4CF00000;
rContents[583] = 32'h18F0F001;
rContents[584] = 32'h820FFFFE;
rContents[585] = 32'h4CF00002;
rContents[586] = 32'h18F0F020;
rContents[587] = 32'h820FFFF7;
rContents[588] = 32'h2F800012;
rContents[589] = 32'h6CF00001;
rContents[590] = 32'h2F010005;
rContents[591] = 32'h6CF00000;
rContents[592] = 32'h4CF00000;
rContents[593] = 32'h18F0F001;
rContents[594] = 32'h820FFFFE;
rContents[595] = 32'h2F800012;
rContents[596] = 32'h6CF00001;
rContents[597] = 32'h2F010005;
rContents[598] = 32'h6CF00000;
rContents[599] = 32'h4CF00000;
rContents[600] = 32'h18F0F001;
rContents[601] = 32'h820FFFFE;
rContents[602] = 32'h4CF00002;
rContents[603] = 32'h41C00000;
rContents[604] = 32'hF0000000;
rContents[605] = 32'h61C00000;
rContents[606] = 32'h61D00000;
rContents[607] = 32'h18111003;
rContents[608] = 32'h41C00000;
rContents[609] = 32'h18011004;
rContents[610] = 32'h2D000020;
rContents[611] = 32'h61D00000;
rContents[612] = 32'hD00FFF95;
rContents[613] = 32'h41D00000;
rContents[614] = 32'h18BFF078;
rContents[615] = 32'h186CC003;
rContents[616] = 32'h103CCF00;
rContents[617] = 32'h61D00000;
rContents[618] = 32'h61C00000;
rContents[619] = 32'hD00FFF77;
rContents[620] = 32'h41C00000;
rContents[621] = 32'h41D00000;
rContents[622] = 32'h41D00000;
rContents[623] = 32'h41C00000;
rContents[624] = 32'hF0000000;
rContents[625] = 32'h61C00000;
rContents[626] = 32'h61D00000;
rContents[627] = 32'h18111003;
rContents[628] = 32'h41C00000;
rContents[629] = 32'h18011004;
rContents[630] = 32'h2D000021;
rContents[631] = 32'h61D00000;
rContents[632] = 32'h61C00000;
rContents[633] = 32'hD00FFF69;
rContents[634] = 32'h41C00000;
rContents[635] = 32'h41D00000;
rContents[636] = 32'h2D000020;
rContents[637] = 32'h61D00000;
rContents[638] = 32'hD00FFF7B;
rContents[639] = 32'h41D00000;
rContents[640] = 32'h183FF080;
rContents[641] = 32'h61D00000;
rContents[642] = 32'h61F00000;
rContents[643] = 32'hD00FFF5F;
rContents[644] = 32'h41F00000;
rContents[645] = 32'h41D00000;
rContents[646] = 32'h2D000020;
rContents[647] = 32'h61D00000;
rContents[648] = 32'hD00FFF71;
rContents[649] = 32'h18F0F080;
rContents[650] = 32'h820FFFFE;
rContents[651] = 32'h41D00000;
rContents[652] = 32'h2D000022;
rContents[653] = 32'h61D00000;
rContents[654] = 32'hD00FFF6B;
rContents[655] = 32'h41D00000;
rContents[656] = 32'h41D00000;
rContents[657] = 32'h41C00000;
rContents[658] = 32'hF0000000;
rContents[659] = 32'h61D00000;
rContents[660] = 32'h2D000021;
rContents[661] = 32'h61D00000;
rContents[662] = 32'h2D0000FF;
rContents[663] = 32'h61D00000;
rContents[664] = 32'hD00FFF4A;
rContents[665] = 32'h41D00000;
rContents[666] = 32'h41D00000;
rContents[667] = 32'h2D000020;
rContents[668] = 32'h61D00000;
rContents[669] = 32'hD00FFF5C;
rContents[670] = 32'h41D00000;
rContents[671] = 32'h183FF080;
rContents[672] = 32'h61D00000;
rContents[673] = 32'h61F00000;
rContents[674] = 32'hD00FFF40;
rContents[675] = 32'h41F00000;
rContents[676] = 32'h41D00000;
rContents[677] = 32'h2D000020;
rContents[678] = 32'h61D00000;
rContents[679] = 32'hD00FFF52;
rContents[680] = 32'h18F0F080;
rContents[681] = 32'h820FFFFE;
rContents[682] = 32'h41D00000;
rContents[683] = 32'h2D000022;
rContents[684] = 32'h61D00000;
rContents[685] = 32'hD00FFF4C;
rContents[686] = 32'h41D00000;
rContents[687] = 32'h41D00000;
rContents[688] = 32'hF0000000;
rContents[689] = 32'h61C00000;
rContents[690] = 32'h61D00000;
rContents[691] = 32'h61E00000;
rContents[692] = 32'h18111004;
rContents[693] = 32'h41C00000;
rContents[694] = 32'h2E000008;
rContents[695] = 32'h18011005;
rContents[696] = 32'h182DCCF0;
rContents[697] = 32'h186CC004;
rContents[698] = 32'h188DD01C;
rContents[699] = 32'h180DD030;
rContents[700] = 32'h18E0D03A;
rContents[701] = 32'h84000002;
rContents[702] = 32'h180DD007;
rContents[703] = 32'h61D00000;
rContents[704] = 32'hD00FFF55;
rContents[705] = 32'hD0000225;
rContents[706] = 32'h41D00000;
rContents[707] = 32'h181EE001;
rContents[708] = 32'h18E0E000;
rContents[709] = 32'h820FFFF3;
rContents[710] = 32'h41E00000;
rContents[711] = 32'h41D00000;
rContents[712] = 32'h41C00000;
rContents[713] = 32'hF0000000;
rContents[714] = 32'h61C00000;
rContents[715] = 32'h61D00000;
rContents[716] = 32'h61E00000;
rContents[717] = 32'h18111004;
rContents[718] = 32'h41D00000;
rContents[719] = 32'h41C00000;
rContents[720] = 32'h18011006;
rContents[721] = 32'h61D00000;
rContents[722] = 32'h61C00000;
rContents[723] = 32'h2C000008;
rContents[724] = 32'h101DCD00;
rContents[725] = 32'h186DD002;
rContents[726] = 32'h41C00000;
rContents[727] = 32'h106CCD00;
rContents[728] = 32'h41D00000;
rContents[729] = 32'h182ECCF0;
rContents[730] = 32'h186CC004;
rContents[731] = 32'h188EE01C;
rContents[732] = 32'h180EE030;
rContents[733] = 32'h18E0E03A;
rContents[734] = 32'h84000002;
rContents[735] = 32'h180EE007;
rContents[736] = 32'h61E00000;
rContents[737] = 32'hD00FFF34;
rContents[738] = 32'hD0000204;
rContents[739] = 32'h41E00000;
rContents[740] = 32'h181DD001;
rContents[741] = 32'h18E0D000;
rContents[742] = 32'h820FFFF3;
rContents[743] = 32'h41E00000;
rContents[744] = 32'h41D00000;
rContents[745] = 32'h41C00000;
rContents[746] = 32'hF0000000;
rContents[747] = 32'h61C00000;
rContents[748] = 32'h61D00000;
rContents[749] = 32'h61E00000;
rContents[750] = 32'h18111004;
rContents[751] = 32'h41D00000;
rContents[752] = 32'h41C00000;
rContents[753] = 32'h18011006;
rContents[754] = 32'h08ED0000;
rContents[755] = 32'h187DD002;
rContents[756] = 32'h100CCD00;
rContents[757] = 32'h4CF00000;
rContents[758] = 32'h2D000003;
rContents[759] = 32'h182EE003;
rContents[760] = 32'h101EDE00;
rContents[761] = 32'h186EE003;
rContents[762] = 32'h10DFFEFF;
rContents[763] = 32'h41E00000;
rContents[764] = 32'h41D00000;
rContents[765] = 32'h41C00000;
rContents[766] = 32'hF0000000;
rContents[767] = 32'h61C00000;
rContents[768] = 32'h61D00000;
rContents[769] = 32'h18111003;
rContents[770] = 32'h2D000000;
rContents[771] = 32'h41C00000;
rContents[772] = 32'h18011004;
rContents[773] = 32'h61C00000;
rContents[774] = 32'h61D00000;
rContents[775] = 32'hD00FFFE4;
rContents[776] = 32'h41D00000;
rContents[777] = 32'h18E0F000;
rContents[778] = 32'h81000007;
rContents[779] = 32'h61F00000;
rContents[780] = 32'hD00FFF09;
rContents[781] = 32'hD00001D9;
rContents[782] = 32'h41F00000;
rContents[783] = 32'h180DD001;
rContents[784] = 32'h800FFFF6;
rContents[785] = 32'h41C00000;
rContents[786] = 32'h41D00000;
rContents[787] = 32'h41C00000;
rContents[788] = 32'hF0000000;
rContents[789] = 32'h61C00000;
rContents[790] = 32'h61D00000;
rContents[791] = 32'h61E00000;
rContents[792] = 32'h18111004;
rContents[793] = 32'h2E000000;
rContents[794] = 32'h41D00000;
rContents[795] = 32'h41C00000;
rContents[796] = 32'h18011006;
rContents[797] = 32'h61C00000;
rContents[798] = 32'h61E00000;
rContents[799] = 32'hD00FFFCC;
rContents[800] = 32'h41E00000;
rContents[801] = 32'h18E0F000;
rContents[802] = 32'h81000009;
rContents[803] = 32'h61F00000;
rContents[804] = 32'hD00FFEF1;
rContents[805] = 32'hD00001C1;
rContents[806] = 32'h41F00000;
rContents[807] = 32'h180EE001;
rContents[808] = 32'h181DD001;
rContents[809] = 32'h18E0D000;
rContents[810] = 32'h820FFFF4;
rContents[811] = 32'h41C00000;
rContents[812] = 32'h41E00000;
rContents[813] = 32'h41D00000;
rContents[814] = 32'h41C00000;
rContents[815] = 32'hF0000000;
rContents[816] = 32'h61C00000;
rContents[817] = 32'h61D00000;
rContents[818] = 32'h61E00000;
rContents[819] = 32'h2C000000;
rContents[820] = 32'h61C00000;
rContents[821] = 32'hD00FFF28;
rContents[822] = 32'h41C00000;
rContents[823] = 32'h2C00000B;
rContents[824] = 32'hD00FFF5B;
rContents[825] = 32'h181CC001;
rContents[826] = 32'h18E0C000;
rContents[827] = 32'h820FFFFD;
rContents[828] = 32'h2C000001;
rContents[829] = 32'h61C00000;
rContents[830] = 32'hD00FFF1F;
rContents[831] = 32'h41C00000;
rContents[832] = 32'h2C000000;
rContents[833] = 32'h61C00000;
rContents[834] = 32'h2C000000;
rContents[835] = 32'h61C00000;
rContents[836] = 32'h2D000001;
rContents[837] = 32'h186DD000;
rContents[838] = 32'h2E000000;
rContents[839] = 32'hD0000084;
rContents[840] = 32'h10E0FD00;
rContents[841] = 32'h81000005;
rContents[842] = 32'h180EE001;
rContents[843] = 32'h18E0E402;
rContents[844] = 32'h8100006E;
rContents[845] = 32'h800FFFFA;
rContents[846] = 32'h41C00000;
rContents[847] = 32'h41C00000;
rContents[848] = 32'h2C000008;
rContents[849] = 32'h61C00000;
rContents[850] = 32'h2C0001AA;
rContents[851] = 32'h61C00000;
rContents[852] = 32'hD0000077;
rContents[853] = 32'h41C00000;
rContents[854] = 32'h41C00000;
rContents[855] = 32'h2D000001;
rContents[856] = 32'h186DD002;
rContents[857] = 32'h10F0FD00;
rContents[858] = 32'h8200000C;
rContents[859] = 32'hD00FFF38;
rContents[860] = 32'hD00FFF37;
rContents[861] = 32'hD00FFF36;
rContents[862] = 32'h18F0F001;
rContents[863] = 32'h8100005D;
rContents[864] = 32'hD00FFF33;
rContents[865] = 32'h18E0F0AA;
rContents[866] = 32'h8200005A;
rContents[867] = 32'h2E000001;
rContents[868] = 32'h186EE001;
rContents[869] = 32'h80000014;
rContents[870] = 32'h2C000037;
rContents[871] = 32'h61C00000;
rContents[872] = 32'h2C000000;
rContents[873] = 32'h61C00000;
rContents[874] = 32'hD0000061;
rContents[875] = 32'h41C00000;
rContents[876] = 32'h41C00000;
rContents[877] = 32'h2C000029;
rContents[878] = 32'h61C00000;
rContents[879] = 32'h2C000000;
rContents[880] = 32'h61C00000;
rContents[881] = 32'hD000005A;
rContents[882] = 32'h41C00000;
rContents[883] = 32'h41C00000;
rContents[884] = 32'h2E000000;
rContents[885] = 32'h10E0FD00;
rContents[886] = 32'h82000003;
rContents[887] = 32'h2E000001;
rContents[888] = 32'h186EE000;
rContents[889] = 32'h2D000000;
rContents[890] = 32'h18F0E003;
rContents[891] = 32'h81000013;
rContents[892] = 32'h2C000037;
rContents[893] = 32'h61C00000;
rContents[894] = 32'h2C000000;
rContents[895] = 32'h61C00000;
rContents[896] = 32'hD000004B;
rContents[897] = 32'h41C00000;
rContents[898] = 32'h41C00000;
rContents[899] = 32'h2C000029;
rContents[900] = 32'h61C00000;
rContents[901] = 32'h2C000000;
rContents[902] = 32'h18F0E002;
rContents[903] = 32'h81000002;
rContents[904] = 32'h2C804000;
rContents[905] = 32'h61C00000;
rContents[906] = 32'hD0000041;
rContents[907] = 32'h41C00000;
rContents[908] = 32'h41C00000;
rContents[909] = 32'h80000008;
rContents[910] = 32'h2C000029;
rContents[911] = 32'h61C00000;
rContents[912] = 32'h2C000000;
rContents[913] = 32'h61C00000;
rContents[914] = 32'hD0000039;
rContents[915] = 32'h41C00000;
rContents[916] = 32'h41C00000;
rContents[917] = 32'h18F0F001;
rContents[918] = 32'h81000005;
rContents[919] = 32'h180DD001;
rContents[920] = 32'h18E0D480;
rContents[921] = 32'h81000023;
rContents[922] = 32'h800FFFE0;
rContents[923] = 32'h18F0E002;
rContents[924] = 32'h81000013;
rContents[925] = 32'h2C00003A;
rContents[926] = 32'h61C00000;
rContents[927] = 32'h2C000000;
rContents[928] = 32'h61C00000;
rContents[929] = 32'hD000002A;
rContents[930] = 32'h41C00000;
rContents[931] = 32'h41C00000;
rContents[932] = 32'h18E0F000;
rContents[933] = 32'h82000017;
rContents[934] = 32'hD00FFEED;
rContents[935] = 32'h18F0F040;
rContents[936] = 32'h81000004;
rContents[937] = 32'h2C000001;
rContents[938] = 32'h186CC002;
rContents[939] = 32'h103EEC00;
rContents[940] = 32'hD00FFEE7;
rContents[941] = 32'hD00FFEE6;
rContents[942] = 32'hD00FFEE5;
rContents[943] = 32'h2C000010;
rContents[944] = 32'h61C00000;
rContents[945] = 32'h2C000200;
rContents[946] = 32'h61C00000;
rContents[947] = 32'hD0000018;
rContents[948] = 32'h41C00000;
rContents[949] = 32'h41C00000;
rContents[950] = 32'h18E0F000;
rContents[951] = 32'h82000005;
rContents[952] = 32'h8000000A;
rContents[953] = 32'hD00001B4;
rContents[954] = 32'h41C00000;
rContents[955] = 32'h41C00000;
rContents[956] = 32'h2C000000;
rContents[957] = 32'h61C00000;
rContents[958] = 32'hD00FFE9F;
rContents[959] = 32'h41C00000;
rContents[960] = 32'h2F0000FF;
rContents[961] = 32'h80000006;
rContents[962] = 32'h2C000000;
rContents[963] = 32'h61C00000;
rContents[964] = 32'hD00FFE99;
rContents[965] = 32'h41C00000;
rContents[966] = 32'h08FE0000;
rContents[967] = 32'h41E00000;
rContents[968] = 32'h41D00000;
rContents[969] = 32'h41C00000;
rContents[970] = 32'hF0000000;
rContents[971] = 32'h61C00000;
rContents[972] = 32'h61D00000;
rContents[973] = 32'h18111003;
rContents[974] = 32'h41D00000;
rContents[975] = 32'h41C00000;
rContents[976] = 32'h18011005;
rContents[977] = 32'hD00FFEC2;
rContents[978] = 32'h183CC040;
rContents[979] = 32'h61C00000;
rContents[980] = 32'hD00FFE9D;
rContents[981] = 32'h41C00000;
rContents[982] = 32'h61C00000;
rContents[983] = 32'h08CD0000;
rContents[984] = 32'h18DDCCFF;
rContents[985] = 32'h61D00000;
rContents[986] = 32'hD00FFE97;
rContents[987] = 32'h41D00000;
rContents[988] = 32'h18DDC8FF;
rContents[989] = 32'h61D00000;
rContents[990] = 32'hD00FFE93;
rContents[991] = 32'h41D00000;
rContents[992] = 32'h18DDC4FF;
rContents[993] = 32'h61D00000;
rContents[994] = 32'hD00FFE8F;
rContents[995] = 32'h41D00000;
rContents[996] = 32'h18DDC0FF;
rContents[997] = 32'h61D00000;
rContents[998] = 32'hD00FFE8B;
rContents[999] = 32'h41D00000;
rContents[1000] = 32'h41C00000;
rContents[1001] = 32'h18E0C040;
rContents[1002] = 32'h82000003;
rContents[1003] = 32'h2D000095;
rContents[1004] = 32'h80000006;
rContents[1005] = 32'h18E0C048;
rContents[1006] = 32'h82000003;
rContents[1007] = 32'h2D000087;
rContents[1008] = 32'h80000002;
rContents[1009] = 32'h2D0000FF;
rContents[1010] = 32'h61D00000;
rContents[1011] = 32'hD00FFE7E;
rContents[1012] = 32'h41D00000;
rContents[1013] = 32'h2D00000A;
rContents[1014] = 32'hD00FFE9D;
rContents[1015] = 32'h18E0F0FF;
rContents[1016] = 32'h82000005;
rContents[1017] = 32'h181DD001;
rContents[1018] = 32'h18E0D000;
rContents[1019] = 32'h81000002;
rContents[1020] = 32'h800FFFFA;
rContents[1021] = 32'h41D00000;
rContents[1022] = 32'h41C00000;
rContents[1023] = 32'hF0000000;
rContents[1024] = 32'h61C00000;
rContents[1025] = 32'h61D00000;
rContents[1026] = 32'h61E00000;
rContents[1027] = 32'h18111004;
rContents[1028] = 32'h41D00000;
rContents[1029] = 32'h41C00000;
rContents[1030] = 32'h18011006;
rContents[1031] = 32'h2F000001;
rContents[1032] = 32'h61F00000;
rContents[1033] = 32'hD00FFE54;
rContents[1034] = 32'h41F00000;
rContents[1035] = 32'h186DD009;
rContents[1036] = 32'h2F000011;
rContents[1037] = 32'h61F00000;
rContents[1038] = 32'h61D00000;
rContents[1039] = 32'hD00FFFBC;
rContents[1040] = 32'h18111002;
rContents[1041] = 32'h18E0F000;
rContents[1042] = 32'h82000023;
rContents[1043] = 32'hD00FFE80;
rContents[1044] = 32'h18E0F0FE;
rContents[1045] = 32'h820FFFFE;
rContents[1046] = 32'h2E000080;
rContents[1047] = 32'h2D000000;
rContents[1048] = 32'hD00FFE7B;
rContents[1049] = 32'h186DF018;
rContents[1050] = 32'hD00FFE79;
rContents[1051] = 32'h186FF010;
rContents[1052] = 32'h103DDF00;
rContents[1053] = 32'hD00FFE76;
rContents[1054] = 32'h186FF008;
rContents[1055] = 32'h103DDF00;
rContents[1056] = 32'hD00FFE73;
rContents[1057] = 32'h103DDF00;
rContents[1058] = 32'h6CD00000;
rContents[1059] = 32'h180CC001;
rContents[1060] = 32'h181EE001;
rContents[1061] = 32'h18E0E000;
rContents[1062] = 32'h820FFFF2;
rContents[1063] = 32'hD00FFE6C;
rContents[1064] = 32'hD00FFE6B;
rContents[1065] = 32'h2F000000;
rContents[1066] = 32'h61F00000;
rContents[1067] = 32'hD00FFE32;
rContents[1068] = 32'h41F00000;
rContents[1069] = 32'hD00FFE66;
rContents[1070] = 32'hD00FFE65;
rContents[1071] = 32'hD00FFE64;
rContents[1072] = 32'hD00FFE63;
rContents[1073] = 32'hD00FFE62;
rContents[1074] = 32'hD00FFE61;
rContents[1075] = 32'h2F000000;
rContents[1076] = 32'h80000009;
rContents[1077] = 32'h61F00000;
rContents[1078] = 32'hD00FFE7B;
rContents[1079] = 32'h41F00000;
rContents[1080] = 32'h2F000000;
rContents[1081] = 32'h61F00000;
rContents[1082] = 32'hD00FFE23;
rContents[1083] = 32'h41F00000;
rContents[1084] = 32'h2F0000FF;
rContents[1085] = 32'h41E00000;
rContents[1086] = 32'h41D00000;
rContents[1087] = 32'h41C00000;
rContents[1088] = 32'hF0000000;
rContents[1089] = 32'h61C00000;
rContents[1090] = 32'h61D00000;
rContents[1091] = 32'h61E00000;
rContents[1092] = 32'h18111004;
rContents[1093] = 32'h41D00000;
rContents[1094] = 32'h41C00000;
rContents[1095] = 32'h18011006;
rContents[1096] = 32'h2F000001;
rContents[1097] = 32'h61F00000;
rContents[1098] = 32'hD00FFE13;
rContents[1099] = 32'h41F00000;
rContents[1100] = 32'h2F000018;
rContents[1101] = 32'h61F00000;
rContents[1102] = 32'h61D00000;
rContents[1103] = 32'hD00FFF7C;
rContents[1104] = 32'h18111002;
rContents[1105] = 32'h18E0F000;
rContents[1106] = 32'h8200002E;
rContents[1107] = 32'h2F0000FE;
rContents[1108] = 32'h61F00000;
rContents[1109] = 32'hD00FFE1C;
rContents[1110] = 32'h41F00000;
rContents[1111] = 32'h2E000080;
rContents[1112] = 32'h4CD00000;
rContents[1113] = 32'h61C00000;
rContents[1114] = 32'h182CDCFF;
rContents[1115] = 32'h188DD018;
rContents[1116] = 32'h61D00000;
rContents[1117] = 32'hD00FFE14;
rContents[1118] = 32'h41D00000;
rContents[1119] = 32'h182CD8FF;
rContents[1120] = 32'h188DD010;
rContents[1121] = 32'h61D00000;
rContents[1122] = 32'hD00FFE0F;
rContents[1123] = 32'h41D00000;
rContents[1124] = 32'h182CD4FF;
rContents[1125] = 32'h188DD008;
rContents[1126] = 32'h61D00000;
rContents[1127] = 32'hD00FFE0A;
rContents[1128] = 32'h41D00000;
rContents[1129] = 32'h182CD0FF;
rContents[1130] = 32'h61D00000;
rContents[1131] = 32'hD00FFE06;
rContents[1132] = 32'h41D00000;
rContents[1133] = 32'h41C00000;
rContents[1134] = 32'h180CC001;
rContents[1135] = 32'h181EE001;
rContents[1136] = 32'h18E0E000;
rContents[1137] = 32'h820FFFE7;
rContents[1138] = 32'h2F0000FF;
rContents[1139] = 32'h61F00000;
rContents[1140] = 32'hD00FFDFD;
rContents[1141] = 32'hD00FFDFC;
rContents[1142] = 32'h41F00000;
rContents[1143] = 32'hD00FFE1C;
rContents[1144] = 32'h18E0F0FF;
rContents[1145] = 32'h820FFFFE;
rContents[1146] = 32'h2F000000;
rContents[1147] = 32'h61F00000;
rContents[1148] = 32'hD00FFDE1;
rContents[1149] = 32'h41F00000;
rContents[1150] = 32'h2F000000;
rContents[1151] = 32'h80000006;
rContents[1152] = 32'h2F000000;
rContents[1153] = 32'h61F00000;
rContents[1154] = 32'hD00FFDDB;
rContents[1155] = 32'h41F00000;
rContents[1156] = 32'h2F0000FF;
rContents[1157] = 32'h41E00000;
rContents[1158] = 32'h41D00000;
rContents[1159] = 32'h41C00000;
rContents[1160] = 32'hF0000000;
rContents[1161] = 32'h61D00000;
rContents[1162] = 32'h2D000030;
rContents[1163] = 32'h61D00000;
rContents[1164] = 32'h2D000000;
rContents[1165] = 32'h61D00000;
rContents[1166] = 32'hD00FFD54;
rContents[1167] = 32'h41D00000;
rContents[1168] = 32'h41D00000;
rContents[1169] = 32'h2D000031;
rContents[1170] = 32'h61D00000;
rContents[1171] = 32'h2D000000;
rContents[1172] = 32'h61D00000;
rContents[1173] = 32'hD00FFD4D;
rContents[1174] = 32'h41D00000;
rContents[1175] = 32'h41D00000;
rContents[1176] = 32'h2D000032;
rContents[1177] = 32'h61D00000;
rContents[1178] = 32'h2D000000;
rContents[1179] = 32'h61D00000;
rContents[1180] = 32'hD00FFD46;
rContents[1181] = 32'h41D00000;
rContents[1182] = 32'h41D00000;
rContents[1183] = 32'hD0000003;
rContents[1184] = 32'h41D00000;
rContents[1185] = 32'hF0000000;
rContents[1186] = 32'h61D00000;
rContents[1187] = 32'h2D000031;
rContents[1188] = 32'h61D00000;
rContents[1189] = 32'h2D000000;
rContents[1190] = 32'h61D00000;
rContents[1191] = 32'hD00FFD3B;
rContents[1192] = 32'h41D00000;
rContents[1193] = 32'h41D00000;
rContents[1194] = 32'h2D000032;
rContents[1195] = 32'h61D00000;
rContents[1196] = 32'h2D000000;
rContents[1197] = 32'h61D00000;
rContents[1198] = 32'hD00FFD34;
rContents[1199] = 32'h41D00000;
rContents[1200] = 32'h41D00000;
rContents[1201] = 32'h2D000033;
rContents[1202] = 32'h61D00000;
rContents[1203] = 32'h2D000000;
rContents[1204] = 32'h61D00000;
rContents[1205] = 32'hD00FFD2D;
rContents[1206] = 32'h41D00000;
rContents[1207] = 32'h41D00000;
rContents[1208] = 32'h2D000031;
rContents[1209] = 32'h61D00000;
rContents[1210] = 32'hD00FFD3F;
rContents[1211] = 32'h41D00000;
rContents[1212] = 32'h180FF001;
rContents[1213] = 32'h61F00000;
rContents[1214] = 32'h2D000031;
rContents[1215] = 32'h61D00000;
rContents[1216] = 32'h61F00000;
rContents[1217] = 32'hD00FFD21;
rContents[1218] = 32'h41F00000;
rContents[1219] = 32'h41D00000;
rContents[1220] = 32'h41F00000;
rContents[1221] = 32'h18E0F050;
rContents[1222] = 32'h820FFFEB;
rContents[1223] = 32'h2D000031;
rContents[1224] = 32'h61D00000;
rContents[1225] = 32'h2D000000;
rContents[1226] = 32'h61D00000;
rContents[1227] = 32'hD00FFD17;
rContents[1228] = 32'h41D00000;
rContents[1229] = 32'h41D00000;
rContents[1230] = 32'h2D000032;
rContents[1231] = 32'h61D00000;
rContents[1232] = 32'hD00FFD29;
rContents[1233] = 32'h41D00000;
rContents[1234] = 32'h180FF001;
rContents[1235] = 32'h61F00000;
rContents[1236] = 32'h2D000032;
rContents[1237] = 32'h61D00000;
rContents[1238] = 32'h61F00000;
rContents[1239] = 32'hD00FFD0B;
rContents[1240] = 32'h41F00000;
rContents[1241] = 32'h41D00000;
rContents[1242] = 32'h41F00000;
rContents[1243] = 32'h18E0F028;
rContents[1244] = 32'h820FFFD5;
rContents[1245] = 32'h2D000032;
rContents[1246] = 32'h61D00000;
rContents[1247] = 32'h2D000000;
rContents[1248] = 32'h61D00000;
rContents[1249] = 32'hD00FFD01;
rContents[1250] = 32'h41D00000;
rContents[1251] = 32'h41D00000;
rContents[1252] = 32'h41D00000;
rContents[1253] = 32'hF0000000;
rContents[1254] = 32'h61C00000;
rContents[1255] = 32'h61D00000;
rContents[1256] = 32'h18111003;
rContents[1257] = 32'h41C00000;
rContents[1258] = 32'h18011004;
rContents[1259] = 32'h18E0C020;
rContents[1260] = 32'h8300001E;
rContents[1261] = 32'h18E0C00D;
rContents[1262] = 32'h82000009;
rContents[1263] = 32'h2D000031;
rContents[1264] = 32'h61D00000;
rContents[1265] = 32'h2D000000;
rContents[1266] = 32'h61D00000;
rContents[1267] = 32'hD00FFCEF;
rContents[1268] = 32'h41D00000;
rContents[1269] = 32'h41D00000;
rContents[1270] = 32'h80000048;
rContents[1271] = 32'h18E0C00A;
rContents[1272] = 32'h82000011;
rContents[1273] = 32'h2D000032;
rContents[1274] = 32'h61D00000;
rContents[1275] = 32'hD00FFCFE;
rContents[1276] = 32'h41D00000;
rContents[1277] = 32'h180FF001;
rContents[1278] = 32'h61F00000;
rContents[1279] = 32'h2D000032;
rContents[1280] = 32'h61D00000;
rContents[1281] = 32'h61F00000;
rContents[1282] = 32'hD00FFCE0;
rContents[1283] = 32'h41F00000;
rContents[1284] = 32'h41D00000;
rContents[1285] = 32'h41F00000;
rContents[1286] = 32'h18E0F028;
rContents[1287] = 32'h81000036;
rContents[1288] = 32'h80000036;
rContents[1289] = 32'h80000035;
rContents[1290] = 32'h183CC4FF;
rContents[1291] = 32'h2D000033;
rContents[1292] = 32'h61D00000;
rContents[1293] = 32'h61C00000;
rContents[1294] = 32'hD00FFCD4;
rContents[1295] = 32'h41C00000;
rContents[1296] = 32'h41D00000;
rContents[1297] = 32'h2D000031;
rContents[1298] = 32'h61D00000;
rContents[1299] = 32'hD00FFCE6;
rContents[1300] = 32'h41D00000;
rContents[1301] = 32'h180FF001;
rContents[1302] = 32'h61F00000;
rContents[1303] = 32'h2D000031;
rContents[1304] = 32'h61D00000;
rContents[1305] = 32'h61F00000;
rContents[1306] = 32'hD00FFCC8;
rContents[1307] = 32'h41F00000;
rContents[1308] = 32'h41D00000;
rContents[1309] = 32'h41F00000;
rContents[1310] = 32'h18E0F050;
rContents[1311] = 32'h8200001F;
rContents[1312] = 32'h2D000031;
rContents[1313] = 32'h61D00000;
rContents[1314] = 32'h2D000000;
rContents[1315] = 32'h61D00000;
rContents[1316] = 32'hD00FFCBE;
rContents[1317] = 32'h41D00000;
rContents[1318] = 32'h41D00000;
rContents[1319] = 32'h2D000032;
rContents[1320] = 32'h61D00000;
rContents[1321] = 32'hD00FFCD0;
rContents[1322] = 32'h41D00000;
rContents[1323] = 32'h180FF001;
rContents[1324] = 32'h61F00000;
rContents[1325] = 32'h2D000032;
rContents[1326] = 32'h61D00000;
rContents[1327] = 32'h61F00000;
rContents[1328] = 32'hD00FFCB2;
rContents[1329] = 32'h41F00000;
rContents[1330] = 32'h41D00000;
rContents[1331] = 32'h41F00000;
rContents[1332] = 32'h18E0F028;
rContents[1333] = 32'h82000009;
rContents[1334] = 32'h2D000032;
rContents[1335] = 32'h61D00000;
rContents[1336] = 32'h2D000000;
rContents[1337] = 32'h61D00000;
rContents[1338] = 32'hD00FFCA8;
rContents[1339] = 32'h41D00000;
rContents[1340] = 32'h41D00000;
rContents[1341] = 32'hD00FFF65;
rContents[1342] = 32'h41D00000;
rContents[1343] = 32'h41C00000;
rContents[1344] = 32'hF0000000;
rContents[1345] = 32'h0A0A416E;
rContents[1346] = 32'h20657272;
rContents[1347] = 32'h6F722068;
rContents[1348] = 32'h6173206F;
rContents[1349] = 32'h63637572;
rContents[1350] = 32'h65642E0A;
rContents[1351] = 32'h00000000;
rContents[1352] = 32'h0A0A4120;
rContents[1353] = 32'h66617461;
rContents[1354] = 32'h6C206572;
rContents[1355] = 32'h726F7220;
rContents[1356] = 32'h68617320;
rContents[1357] = 32'h6F636375;
rContents[1358] = 32'h7265642E;
rContents[1359] = 32'h0A000000;
rContents[1360] = 32'h43616C6C;
rContents[1361] = 32'h65642061;
rContents[1362] = 32'h74200000;
rContents[1363] = 32'h53746163;
rContents[1364] = 32'h6B747261;
rContents[1365] = 32'h63652028;
rContents[1366] = 32'h746F7020;
rContents[1367] = 32'h3136293A;
rContents[1368] = 32'h0A000000;
rContents[1369] = 32'h52656769;
rContents[1370] = 32'h73746572;
rContents[1371] = 32'h733A0A00;
rContents[1372] = 32'h52657375;
rContents[1373] = 32'h6D696E67;
rContents[1374] = 32'h2E0A0A00;
rContents[1375] = 32'h48616C74;
rContents[1376] = 32'h696E672E;
rContents[1377] = 32'h0A0A0000;
rContents[1378] = 32'h80000001;
rContents[1379] = 32'h2F000548;
rContents[1380] = 32'h61F00000;
rContents[1381] = 32'hD00FFD9A;
rContents[1382] = 32'h41F00000;
rContents[1383] = 32'h2F000550;
rContents[1384] = 32'h61F00000;
rContents[1385] = 32'hD00FFD96;
rContents[1386] = 32'h41F00000;
rContents[1387] = 32'hD00FFD46;
rContents[1388] = 32'h04200000;
rContents[1389] = 32'h61F00000;
rContents[1390] = 32'h2F000550;
rContents[1391] = 32'h61F00000;
rContents[1392] = 32'hD00FFD8F;
rContents[1393] = 32'h41F00000;
rContents[1394] = 32'h2F0000F0;
rContents[1395] = 32'h181FF001;
rContents[1396] = 32'h18E0F000;
rContents[1397] = 32'h820FFFFE;
rContents[1398] = 32'h18111001;
rContents[1399] = 32'hD00FFD3A;
rContents[1400] = 32'h18011001;
rContents[1401] = 32'h2F00000A;
rContents[1402] = 32'h61F00000;
rContents[1403] = 32'hD0000013;
rContents[1404] = 32'h41F00000;
rContents[1405] = 32'h2F00000D;
rContents[1406] = 32'h61F00000;
rContents[1407] = 32'hD000000F;
rContents[1408] = 32'h41F00000;
rContents[1409] = 32'h41F00000;
rContents[1410] = 32'hF0000000;
rContents[1411] = 32'hF0000000;
rContents[1412] = 32'hF0000000;
rContents[1413] = 32'h4C656D6F;
rContents[1414] = 32'h6E207630;
rContents[1415] = 32'h2E32202D;
rContents[1416] = 32'h20666F72;
rContents[1417] = 32'h20657052;
rContents[1418] = 32'h49534320;
rContents[1419] = 32'h76352073;
rContents[1420] = 32'h79737465;
rContents[1421] = 32'h6D730000;
rContents[1422] = 32'h18111001;
rContents[1423] = 32'h41F00000;
rContents[1424] = 32'h18011002;
rContents[1425] = 32'h61F00000;
rContents[1426] = 32'hD00FFC83;
rContents[1427] = 32'hD00FFF53;
rContents[1428] = 32'h41F00000;
rContents[1429] = 32'hF0000000;
rContents[1430] = 32'h800FFC7F;
rContents[1431] = 32'h800FFF4F;
rContents[1432] = 32'h800FFC99;
rContents[1433] = 32'h800FFD18;
rContents[1434] = 32'h800FFD65;
rContents[1435] = 32'h800FFFC8;
rContents[1436] = 32'h210017FF;
rContents[1437] = 32'h28000585;
rContents[1438] = 32'h61800000;
rContents[1439] = 32'hD00FFFFB;
rContents[1440] = 32'h41800000;
rContents[1441] = 32'h26001000;
rContents[1442] = 32'h29000000;
rContents[1443] = 32'h2800000A;
rContents[1444] = 32'h61800000;
rContents[1445] = 32'hD00FFFE9;
rContents[1446] = 32'h41800000;
rContents[1447] = 32'h2800000D;
rContents[1448] = 32'h61800000;
rContents[1449] = 32'hD00FFFE5;
rContents[1450] = 32'h41800000;
rContents[1451] = 32'h2800003E;
rContents[1452] = 32'h61800000;
rContents[1453] = 32'hD00FFFE1;
rContents[1454] = 32'h41800000;
rContents[1455] = 32'hD00FFFE9;
rContents[1456] = 32'h18E0F008;
rContents[1457] = 32'h8200000E;
rContents[1458] = 32'h18E06000;
rContents[1459] = 32'h82000002;
rContents[1460] = 32'h800FFFFB;
rContents[1461] = 32'h18166002;
rContents[1462] = 32'h18199001;
rContents[1463] = 32'h46F00000;
rContents[1464] = 32'h61F00000;
rContents[1465] = 32'hD00FFFD5;
rContents[1466] = 32'h41F00000;
rContents[1467] = 32'h18066001;
rContents[1468] = 32'h2F000000;
rContents[1469] = 32'h66F00000;
rContents[1470] = 32'h800FFFF1;
rContents[1471] = 32'h18E0F00D;
rContents[1472] = 32'h82000003;
rContents[1473] = 32'h66F00000;
rContents[1474] = 32'h8000000A;
rContents[1475] = 32'h18F09180;
rContents[1476] = 32'h820FFFEB;
rContents[1477] = 32'h61F00000;
rContents[1478] = 32'hD00FFFC8;
rContents[1479] = 32'h41F00000;
rContents[1480] = 32'h66F00000;
rContents[1481] = 32'h18066001;
rContents[1482] = 32'h18099001;
rContents[1483] = 32'h800FFFE4;
rContents[1484] = 32'h26001000;
rContents[1485] = 32'h27000000;
rContents[1486] = 32'h46900000;
rContents[1487] = 32'h18E0900D;
rContents[1488] = 32'h82000005;
rContents[1489] = 32'h18E0703A;
rContents[1490] = 32'h82000002;
rContents[1491] = 32'h41800000;
rContents[1492] = 32'h800FFFCD;
rContents[1493] = 32'h18E09052;
rContents[1494] = 32'h8200000C;
rContents[1495] = 32'h2800000A;
rContents[1496] = 32'h61800000;
rContents[1497] = 32'hD00FFFB5;
rContents[1498] = 32'h41800000;
rContents[1499] = 32'h2800000D;
rContents[1500] = 32'h61800000;
rContents[1501] = 32'hD00FFFB1;
rContents[1502] = 32'h41800000;
rContents[1503] = 32'hD0400000;
rContents[1504] = 32'h18066001;
rContents[1505] = 32'h800FFFED;
rContents[1506] = 32'h18E0903A;
rContents[1507] = 32'h82000005;
rContents[1508] = 32'h2700003A;
rContents[1509] = 32'h61400000;
rContents[1510] = 32'h18066001;
rContents[1511] = 32'h800FFFE7;
rContents[1512] = 32'h18E0902E;
rContents[1513] = 32'h82000007;
rContents[1514] = 32'h18E0703A;
rContents[1515] = 32'h82000002;
rContents[1516] = 32'h41800000;
rContents[1517] = 32'h2700002E;
rContents[1518] = 32'h18066001;
rContents[1519] = 32'h800FFFDF;
rContents[1520] = 32'h18E09020;
rContents[1521] = 32'h82000003;
rContents[1522] = 32'h18066001;
rContents[1523] = 32'h800FFFDB;
rContents[1524] = 32'h25000000;
rContents[1525] = 32'h46900000;
rContents[1526] = 32'h18199030;
rContents[1527] = 32'h18E0900A;
rContents[1528] = 32'h84000007;
rContents[1529] = 32'h18199007;
rContents[1530] = 32'h18E0900A;
rContents[1531] = 32'h84000008;
rContents[1532] = 32'h18E09010;
rContents[1533] = 32'h84000002;
rContents[1534] = 32'h80000005;
rContents[1535] = 32'h18655004;
rContents[1536] = 32'h10355900;
rContents[1537] = 32'h18066001;
rContents[1538] = 32'h800FFFF3;
rContents[1539] = 32'h46900000;
rContents[1540] = 32'h18E0703A;
rContents[1541] = 32'h82000004;
rContents[1542] = 32'h64500000;
rContents[1543] = 32'h18044001;
rContents[1544] = 32'h800FFFC6;
rContents[1545] = 32'h61400000;
rContents[1546] = 32'h08450000;
rContents[1547] = 32'h18E0902E;
rContents[1548] = 32'h82000003;
rContents[1549] = 32'h41800000;
rContents[1550] = 32'h800FFFC0;
rContents[1551] = 32'h18E07000;
rContents[1552] = 32'h82000016;
rContents[1553] = 32'h41800000;
rContents[1554] = 32'h2800000A;
rContents[1555] = 32'h61800000;
rContents[1556] = 32'hD00FFF7A;
rContents[1557] = 32'h41800000;
rContents[1558] = 32'h2800000D;
rContents[1559] = 32'h61800000;
rContents[1560] = 32'hD00FFF76;
rContents[1561] = 32'h41800000;
rContents[1562] = 32'h61400000;
rContents[1563] = 32'hD00FFC96;
rContents[1564] = 32'h41400000;
rContents[1565] = 32'h2800003A;
rContents[1566] = 32'h61800000;
rContents[1567] = 32'hD00FFF6F;
rContents[1568] = 32'h41800000;
rContents[1569] = 32'h44800000;
rContents[1570] = 32'h61800000;
rContents[1571] = 32'hD00FFF76;
rContents[1572] = 32'h41800000;
rContents[1573] = 32'h800FFFA9;
rContents[1574] = 32'h18E0702E;
rContents[1575] = 32'hD20FFF74;
rContents[1576] = 32'h08840000;
rContents[1577] = 32'h41400000;
rContents[1578] = 32'h10E08400;
rContents[1579] = 32'h8B000002;
rContents[1580] = 32'h08840000;
rContents[1581] = 32'h101A8400;
rContents[1582] = 32'h180AA001;
rContents[1583] = 32'h61400000;
rContents[1584] = 32'h2800000A;
rContents[1585] = 32'h61800000;
rContents[1586] = 32'hD00FFF65;
rContents[1587] = 32'h41800000;
rContents[1588] = 32'h2800000A;
rContents[1589] = 32'h61800000;
rContents[1590] = 32'hD00FFF60;
rContents[1591] = 32'h41800000;
rContents[1592] = 32'h2800000D;
rContents[1593] = 32'h61800000;
rContents[1594] = 32'hD00FFF54;
rContents[1595] = 32'h41800000;
rContents[1596] = 32'h61400000;
rContents[1597] = 32'hD00FFC74;
rContents[1598] = 32'h41400000;
rContents[1599] = 32'h2800003A;
rContents[1600] = 32'h61800000;
rContents[1601] = 32'hD00FFF4D;
rContents[1602] = 32'h41800000;
rContents[1603] = 32'h18E0A008;
rContents[1604] = 32'h83000003;
rContents[1605] = 32'h08BA0000;
rContents[1606] = 32'h80000002;
rContents[1607] = 32'h2B000008;
rContents[1608] = 32'h101AAB00;
rContents[1609] = 32'h80000005;
rContents[1610] = 32'h28000020;
rContents[1611] = 32'h61800000;
rContents[1612] = 32'hD00FFF42;
rContents[1613] = 32'h41800000;
rContents[1614] = 32'h44800000;
rContents[1615] = 32'h61800000;
rContents[1616] = 32'hD00FFF49;
rContents[1617] = 32'h41800000;
rContents[1618] = 32'h18044001;
rContents[1619] = 32'h181BB001;
rContents[1620] = 32'h18E0B000;
rContents[1621] = 32'h820FFFF5;
rContents[1622] = 32'h18E0A000;
rContents[1623] = 32'h820FFFDD;
rContents[1624] = 32'h41400000;
rContents[1625] = 32'h27000000;
rContents[1626] = 32'h800FFF74;
    end

endmodule

/*  Program 1 - square wave generator over GPIO
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808000;
        rContents[8] = 32'h3500FFFF;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25000000;
        rContents[17] = 32'h08650000;
        rContents[18] = 32'h36808002;
        rContents[19] = 32'h64600001;
        rContents[20] = 32'h27010005;
        rContents[21] = 32'h64700000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h04000000;
        rContents[26] = 32'h18B5580F;
        rContents[27] = 32'h18055001;
        rContents[28] = 32'h800FFFF5;
        rContents[29] = 32'h0;
        rContents[30] = 32'h0;
        rContents[31] = 32'h0;
        rContents[32] = 32'h0;
        rContents[33] = 32'h0;
        rContents[34] = 32'h0;
        rContents[35] = 32'h0; */
        
/*  Program 2 - print some 'H's over the serial link
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808101;
        rContents[8] = 32'h35000048;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25808100;
        rContents[17] = 32'h35000080;
        rContents[18] = 32'h64500001;
        rContents[19] = 32'h27010005;
        rContents[20] = 32'h64700000;
        rContents[21] = 32'h04000000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h800FFFED; */
