module epRISC_embeddedROM(iClk, iAddr, oData, iEnable);

    input iClk, iEnable;
    input [11:0] iAddr;
    output wire [31:0] oData;
    
    reg [31:0] rDataOut, rContents[0:4095];
    
    assign oData = (iEnable) ? rDataOut : 32'bz;
    
    always @(posedge iClk) begin
        rDataOut = rContents[iAddr];
    end
    
    initial begin
rContents[0] = 32'h21001100;
rContents[1] = 32'h23000000;
rContents[2] = 32'hD00000FC;
rContents[3] = 32'h24007FFF;
rContents[4] = 32'h61400000;
rContents[5] = 32'h24000000;
rContents[6] = 32'h61400000;
rContents[7] = 32'hD0000104;
rContents[8] = 32'h41400000;
rContents[9] = 32'h41400000;
rContents[10] = 32'hD0000364;
rContents[11] = 32'h24000048;
rContents[12] = 32'h61400000;
rContents[13] = 32'hD00001FB;
rContents[14] = 32'h41400000;
rContents[15] = 32'h240000CA;
rContents[16] = 32'h61400000;
rContents[17] = 32'hD00001F7;
rContents[18] = 32'h41400000;
rContents[19] = 32'h240000EC;
rContents[20] = 32'h61400000;
rContents[21] = 32'hD00001F3;
rContents[22] = 32'h41400000;
rContents[23] = 32'h24000041;
rContents[24] = 32'h61400000;
rContents[25] = 32'hD0000181;
rContents[26] = 32'h41400000;
rContents[27] = 32'h24000059;
rContents[28] = 32'h61400000;
rContents[29] = 32'hD00001EB;
rContents[30] = 32'h41400000;
rContents[31] = 32'hD00001FF;
rContents[32] = 32'h24000078;
rContents[33] = 32'h18E0F0FF;
rContents[34] = 32'h81000002;
rContents[35] = 32'h2400006F;
rContents[36] = 32'h61400000;
rContents[37] = 32'hD00001E3;
rContents[38] = 32'h41400000;
rContents[39] = 32'h24003000;
rContents[40] = 32'h61400000;
rContents[41] = 32'h24000000;
rContents[42] = 32'h61400000;
rContents[43] = 32'hD00002C3;
rContents[44] = 32'h41400000;
rContents[45] = 32'h41400000;
rContents[46] = 32'h240000F8;
rContents[47] = 32'h61400000;
rContents[48] = 32'hD00001D8;
rContents[49] = 32'h41400000;
rContents[50] = 32'h8000044D;
rContents[51] = 32'h43F01FF0;
rContents[52] = 32'h61F00000;
rContents[53] = 32'hD0000165;
rContents[54] = 32'h63F01FF1;
rContents[55] = 32'h41F00000;
rContents[56] = 32'hF0000000;
rContents[57] = 32'hD0000183;
rContents[58] = 32'h63F01FF1;
rContents[59] = 32'hF0000000;
rContents[60] = 32'h43F01FF2;
rContents[61] = 32'h61F00000;
rContents[62] = 32'h43F01FF3;
rContents[63] = 32'h61F00000;
rContents[64] = 32'hD0000279;
rContents[65] = 32'h63F01FF4;
rContents[66] = 32'h41F00000;
rContents[67] = 32'h41F00000;
rContents[68] = 32'hF0000000;
rContents[69] = 32'hD00001D9;
rContents[70] = 32'h63F01FF5;
rContents[71] = 32'hF0000000;
rContents[72] = 32'h65705249;
rContents[73] = 32'h53432042;
rContents[74] = 32'h6F6F746C;
rContents[75] = 32'h6F616465;
rContents[76] = 32'h72207633;
rContents[77] = 32'h2E320A0D;
rContents[78] = 32'h636F7079;
rContents[79] = 32'h72696768;
rContents[80] = 32'h74203230;
rContents[81] = 32'h31352D32;
rContents[82] = 32'h30313720;
rContents[83] = 32'h50726F70;
rContents[84] = 32'h6F727469;
rContents[85] = 32'h6F6E616C;
rContents[86] = 32'h204C6162;
rContents[87] = 32'h730A0D0A;
rContents[88] = 32'h0D000000;
rContents[89] = 32'h41747465;
rContents[90] = 32'h6D707469;
rContents[91] = 32'h6E672074;
rContents[92] = 32'h6F206D6F;
rContents[93] = 32'h756E7420;
rContents[94] = 32'h53442063;
rContents[95] = 32'h61726420;
rContents[96] = 32'h696E2073;
rContents[97] = 32'h6C6F7420;
rContents[98] = 32'h412E2E2E;
rContents[99] = 32'h0A0D0000;
rContents[100] = 32'h41747465;
rContents[101] = 32'h6D707469;
rContents[102] = 32'h6E672074;
rContents[103] = 32'h6F206D6F;
rContents[104] = 32'h756E7420;
rContents[105] = 32'h53442063;
rContents[106] = 32'h61726420;
rContents[107] = 32'h696E2073;
rContents[108] = 32'h6C6F7420;
rContents[109] = 32'h422E2E2E;
rContents[110] = 32'h0A0D0000;
rContents[111] = 32'h20205344;
rContents[112] = 32'h20636172;
rContents[113] = 32'h64206D6F;
rContents[114] = 32'h756E7465;
rContents[115] = 32'h64207375;
rContents[116] = 32'h63636573;
rContents[117] = 32'h7366756C;
rContents[118] = 32'h6C792E0A;
rContents[119] = 32'h0D0A0D00;
rContents[120] = 32'h20204572;
rContents[121] = 32'h726F7220;
rContents[122] = 32'h6D6F756E;
rContents[123] = 32'h74696E67;
rContents[124] = 32'h20534420;
rContents[125] = 32'h63617264;
rContents[126] = 32'h2E0A0D0A;
rContents[127] = 32'h0D000000;
rContents[128] = 32'h46657463;
rContents[129] = 32'h68696E67;
rContents[130] = 32'h20646973;
rContents[131] = 32'h6B20696E;
rContents[132] = 32'h666F2E2E;
rContents[133] = 32'h2E0A0D00;
rContents[134] = 32'h20204469;
rContents[135] = 32'h736B2061;
rContents[136] = 32'h70706561;
rContents[137] = 32'h72732074;
rContents[138] = 32'h6F206265;
rContents[139] = 32'h20636F72;
rContents[140] = 32'h72757074;
rContents[141] = 32'h2E0A0D0A;
rContents[142] = 32'h0D000000;
rContents[143] = 32'h2020466F;
rContents[144] = 32'h756E6420;
rContents[145] = 32'h6469736B;
rContents[146] = 32'h20270000;
rContents[147] = 32'h27206174;
rContents[148] = 32'h20626C6F;
rContents[149] = 32'h636B2030;
rContents[150] = 32'h2E0A0D00;
rContents[151] = 32'h20204469;
rContents[152] = 32'h736B2061;
rContents[153] = 32'h70706561;
rContents[154] = 32'h72732074;
rContents[155] = 32'h6F206265;
rContents[156] = 32'h20656D70;
rContents[157] = 32'h74792E0A;
rContents[158] = 32'h0D0A0D00;
rContents[159] = 32'h2020466F;
rContents[160] = 32'h756E6420;
rContents[161] = 32'h00000000;
rContents[162] = 32'h20656E74;
rContents[163] = 32'h72696573;
rContents[164] = 32'h206F6E20;
rContents[165] = 32'h6469736B;
rContents[166] = 32'h2E0A0D0A;
rContents[167] = 32'h0D000000;
rContents[168] = 32'h41766169;
rContents[169] = 32'h6C61626C;
rContents[170] = 32'h6520656E;
rContents[171] = 32'h74726965;
rContents[172] = 32'h733A0A0D;
rContents[173] = 32'h00000000;
rContents[174] = 32'h2020456E;
rContents[175] = 32'h74727920;
rContents[176] = 32'h27000000;
rContents[177] = 32'h273A2073;
rContents[178] = 32'h74617274;
rContents[179] = 32'h20000000;
rContents[180] = 32'h2C206C65;
rContents[181] = 32'h6E677468;
rContents[182] = 32'h20000000;
rContents[183] = 32'h2C206C6F;
rContents[184] = 32'h6164200A;
rContents[185] = 32'h0D000000;
rContents[186] = 32'h53656C65;
rContents[187] = 32'h63742061;
rContents[188] = 32'h6E20656E;
rContents[189] = 32'h74727920;
rContents[190] = 32'h746F2065;
rContents[191] = 32'h78656375;
rContents[192] = 32'h74652C20;
rContents[193] = 32'h6F722074;
rContents[194] = 32'h79706520;
rContents[195] = 32'h276D2720;
rContents[196] = 32'h746F2065;
rContents[197] = 32'h6E746572;
rContents[198] = 32'h20746865;
rContents[199] = 32'h206D6F6E;
rContents[200] = 32'h69746F72;
rContents[201] = 32'h3A000000;
rContents[202] = 32'h53746172;
rContents[203] = 32'h74696E67;
rContents[204] = 32'h20504F53;
rContents[205] = 32'h54732E2E;
rContents[206] = 32'h2E0A0D00;
rContents[207] = 32'h20204D65;
rContents[208] = 32'h6D6F7279;
rContents[209] = 32'h20202020;
rContents[210] = 32'h20202020;
rContents[211] = 32'h20200000;
rContents[212] = 32'h20205541;
rContents[213] = 32'h52542020;
rContents[214] = 32'h20202020;
rContents[215] = 32'h20202020;
rContents[216] = 32'h20200000;
rContents[217] = 32'h20205350;
rContents[218] = 32'h49202020;
rContents[219] = 32'h20202020;
rContents[220] = 32'h20202020;
rContents[221] = 32'h20200000;
rContents[222] = 32'h20207379;
rContents[223] = 32'h73582042;
rContents[224] = 32'h75732020;
rContents[225] = 32'h20202020;
rContents[226] = 32'h20200000;
rContents[227] = 32'h2020492F;
rContents[228] = 32'h4F20436F;
rContents[229] = 32'h6E74726F;
rContents[230] = 32'h6C6C6572;
rContents[231] = 32'h20200000;
rContents[232] = 32'h4F4B0A0D;
rContents[233] = 32'h00000000;
rContents[234] = 32'h4641494C;
rContents[235] = 32'h0A0D0000;
rContents[236] = 32'h504F5354;
rContents[237] = 32'h20737563;
rContents[238] = 32'h63657373;
rContents[239] = 32'h66756C2E;
rContents[240] = 32'h0A0D0A0D;
rContents[241] = 32'h00000000;
rContents[242] = 32'h504F5354;
rContents[243] = 32'h20756E73;
rContents[244] = 32'h75636365;
rContents[245] = 32'h73736675;
rContents[246] = 32'h6C2E0A0D;
rContents[247] = 32'h0A0D0000;
rContents[248] = 32'h456E7465;
rContents[249] = 32'h72696E67;
rContents[250] = 32'h206D6F6E;
rContents[251] = 32'h69746F72;
rContents[252] = 32'h2E2E2E0A;
rContents[253] = 32'h0D0A0D00;
rContents[254] = 32'h61C00000;
rContents[255] = 32'h2C002000;
rContents[256] = 32'h2F010001;
rContents[257] = 32'h6CF00000;
rContents[258] = 32'h04000000;
rContents[259] = 32'h04000000;
rContents[260] = 32'h04000000;
rContents[261] = 32'h04000000;
rContents[262] = 32'h4CF00000;
rContents[263] = 32'h18F0F001;
rContents[264] = 32'h820FFFFE;
rContents[265] = 32'h41C00000;
rContents[266] = 32'hF0000000;
rContents[267] = 32'h61E00000;
rContents[268] = 32'h61D00000;
rContents[269] = 32'h61C00000;
rContents[270] = 32'h18111004;
rContents[271] = 32'h2C002000;
rContents[272] = 32'h41D00000;
rContents[273] = 32'h41E00000;
rContents[274] = 32'h18011006;
rContents[275] = 32'h2F600008;
rContents[276] = 32'h103FFE00;
rContents[277] = 32'h186FF010;
rContents[278] = 32'h103FFD00;
rContents[279] = 32'h6CF00001;
rContents[280] = 32'h2F010005;
rContents[281] = 32'h6CF00000;
rContents[282] = 32'h4CF00000;
rContents[283] = 32'h18F0F001;
rContents[284] = 32'h820FFFFE;
rContents[285] = 32'h4CF00002;
rContents[286] = 32'h41C00000;
rContents[287] = 32'h41D00000;
rContents[288] = 32'h41E00000;
rContents[289] = 32'hF0000000;
rContents[290] = 32'h61E00000;
rContents[291] = 32'h61C00000;
rContents[292] = 32'h18111003;
rContents[293] = 32'h2C002000;
rContents[294] = 32'h41E00000;
rContents[295] = 32'h18011004;
rContents[296] = 32'h2F600000;
rContents[297] = 32'h103FFE00;
rContents[298] = 32'h186FF010;
rContents[299] = 32'h6CF00001;
rContents[300] = 32'h2F010005;
rContents[301] = 32'h6CF00000;
rContents[302] = 32'h4CF00000;
rContents[303] = 32'h18F0F001;
rContents[304] = 32'h820FFFFE;
rContents[305] = 32'h2F600000;
rContents[306] = 32'h103FFE00;
rContents[307] = 32'h186FF010;
rContents[308] = 32'h6CF00001;
rContents[309] = 32'h2F010005;
rContents[310] = 32'h6CF00000;
rContents[311] = 32'h4CF00000;
rContents[312] = 32'h18F0F001;
rContents[313] = 32'h820FFFFE;
rContents[314] = 32'h4CF00002;
rContents[315] = 32'h41C00000;
rContents[316] = 32'h41E00000;
rContents[317] = 32'hF0000000;
rContents[318] = 32'h61D00000;
rContents[319] = 32'h61C00000;
rContents[320] = 32'h18111003;
rContents[321] = 32'h2C002000;
rContents[322] = 32'h41D00000;
rContents[323] = 32'h18011004;
rContents[324] = 32'h2F000011;
rContents[325] = 32'h61F00000;
rContents[326] = 32'h61D00000;
rContents[327] = 32'hD00FFFC4;
rContents[328] = 32'h41D00000;
rContents[329] = 32'h41F00000;
rContents[330] = 32'h2F000010;
rContents[331] = 32'h61F00000;
rContents[332] = 32'h2F000080;
rContents[333] = 32'h61F00000;
rContents[334] = 32'hD00FFFBD;
rContents[335] = 32'h41D00000;
rContents[336] = 32'h41F00000;
rContents[337] = 32'h2F000010;
rContents[338] = 32'h61F00000;
rContents[339] = 32'hD00FFFCF;
rContents[340] = 32'h18F0F080;
rContents[341] = 32'h820FFFFE;
rContents[342] = 32'h41F00000;
rContents[343] = 32'h41C00000;
rContents[344] = 32'h41D00000;
rContents[345] = 32'hF0000000;
rContents[346] = 32'h61C00000;
rContents[347] = 32'h2C002000;
rContents[348] = 32'h2F808010;
rContents[349] = 32'h3F000020;
rContents[350] = 32'h6CF00001;
rContents[351] = 32'h2F010005;
rContents[352] = 32'h6CF00000;
rContents[353] = 32'h4CF00000;
rContents[354] = 32'h18F0F001;
rContents[355] = 32'h820FFFFE;
rContents[356] = 32'h2F800010;
rContents[357] = 32'h6CF00001;
rContents[358] = 32'h2F010005;
rContents[359] = 32'h6CF00000;
rContents[360] = 32'h4CF00000;
rContents[361] = 32'h18F0F001;
rContents[362] = 32'h820FFFFE;
rContents[363] = 32'h2F800010;
rContents[364] = 32'h6CF00001;
rContents[365] = 32'h2F010005;
rContents[366] = 32'h6CF00000;
rContents[367] = 32'h4CF00000;
rContents[368] = 32'h18F0F001;
rContents[369] = 32'h820FFFFE;
rContents[370] = 32'h4CF00002;
rContents[371] = 32'h18F0F020;
rContents[372] = 32'h820FFFF7;
rContents[373] = 32'h2F800012;
rContents[374] = 32'h6CF00001;
rContents[375] = 32'h2F010005;
rContents[376] = 32'h6CF00000;
rContents[377] = 32'h4CF00000;
rContents[378] = 32'h18F0F001;
rContents[379] = 32'h820FFFFE;
rContents[380] = 32'h2F800012;
rContents[381] = 32'h6CF00001;
rContents[382] = 32'h2F010005;
rContents[383] = 32'h6CF00000;
rContents[384] = 32'h4CF00000;
rContents[385] = 32'h18F0F001;
rContents[386] = 32'h820FFFFE;
rContents[387] = 32'h4CF00002;
rContents[388] = 32'h41C00000;
rContents[389] = 32'hF0000000;
rContents[390] = 32'h61C00000;
rContents[391] = 32'h61D00000;
rContents[392] = 32'h18111003;
rContents[393] = 32'h41C00000;
rContents[394] = 32'h18011004;
rContents[395] = 32'h2D000020;
rContents[396] = 32'h61D00000;
rContents[397] = 32'hD00FFF95;
rContents[398] = 32'h41D00000;
rContents[399] = 32'h18BFF078;
rContents[400] = 32'h186CC003;
rContents[401] = 32'h103CCF00;
rContents[402] = 32'h61D00000;
rContents[403] = 32'h61C00000;
rContents[404] = 32'hD00FFF77;
rContents[405] = 32'h41C00000;
rContents[406] = 32'h41D00000;
rContents[407] = 32'h41D00000;
rContents[408] = 32'h41C00000;
rContents[409] = 32'hF0000000;
rContents[410] = 32'h61C00000;
rContents[411] = 32'h61D00000;
rContents[412] = 32'h18111003;
rContents[413] = 32'h41C00000;
rContents[414] = 32'h18011004;
rContents[415] = 32'h2D000021;
rContents[416] = 32'h61D00000;
rContents[417] = 32'h61C00000;
rContents[418] = 32'hD00FFF69;
rContents[419] = 32'h41C00000;
rContents[420] = 32'h41D00000;
rContents[421] = 32'h2D000020;
rContents[422] = 32'h61D00000;
rContents[423] = 32'hD00FFF7B;
rContents[424] = 32'h41D00000;
rContents[425] = 32'h183FF080;
rContents[426] = 32'h61D00000;
rContents[427] = 32'h61F00000;
rContents[428] = 32'hD00FFF5F;
rContents[429] = 32'h41F00000;
rContents[430] = 32'h41D00000;
rContents[431] = 32'h2D000020;
rContents[432] = 32'h61D00000;
rContents[433] = 32'hD00FFF71;
rContents[434] = 32'h18F0F080;
rContents[435] = 32'h820FFFFE;
rContents[436] = 32'h41D00000;
rContents[437] = 32'h2D000022;
rContents[438] = 32'h61D00000;
rContents[439] = 32'hD00FFF6B;
rContents[440] = 32'h41D00000;
rContents[441] = 32'h41D00000;
rContents[442] = 32'h41C00000;
rContents[443] = 32'hF0000000;
rContents[444] = 32'h61D00000;
rContents[445] = 32'h2D000021;
rContents[446] = 32'h61D00000;
rContents[447] = 32'h2D0000FF;
rContents[448] = 32'h61D00000;
rContents[449] = 32'hD00FFF4A;
rContents[450] = 32'h41D00000;
rContents[451] = 32'h41D00000;
rContents[452] = 32'h2D000020;
rContents[453] = 32'h61D00000;
rContents[454] = 32'hD00FFF5C;
rContents[455] = 32'h41D00000;
rContents[456] = 32'h183FF080;
rContents[457] = 32'h61D00000;
rContents[458] = 32'h61F00000;
rContents[459] = 32'hD00FFF40;
rContents[460] = 32'h41F00000;
rContents[461] = 32'h41D00000;
rContents[462] = 32'h2D000020;
rContents[463] = 32'h61D00000;
rContents[464] = 32'hD00FFF52;
rContents[465] = 32'h18F0F080;
rContents[466] = 32'h820FFFFE;
rContents[467] = 32'h41D00000;
rContents[468] = 32'h2D000022;
rContents[469] = 32'h61D00000;
rContents[470] = 32'hD00FFF4C;
rContents[471] = 32'h41D00000;
rContents[472] = 32'h41D00000;
rContents[473] = 32'hF0000000;
rContents[474] = 32'h61C00000;
rContents[475] = 32'h61D00000;
rContents[476] = 32'h61E00000;
rContents[477] = 32'h18111004;
rContents[478] = 32'h41C00000;
rContents[479] = 32'h2E000008;
rContents[480] = 32'h18011005;
rContents[481] = 32'h182DCCF0;
rContents[482] = 32'h186CC004;
rContents[483] = 32'h188DD01C;
rContents[484] = 32'h180DD030;
rContents[485] = 32'h18E0D03A;
rContents[486] = 32'h84000003;
rContents[487] = 32'h18B22008;
rContents[488] = 32'h180DD007;
rContents[489] = 32'h61D00000;
rContents[490] = 32'hD00FFF54;
rContents[491] = 32'hD00001E0;
rContents[492] = 32'h41D00000;
rContents[493] = 32'h181EE001;
rContents[494] = 32'h18E0E000;
rContents[495] = 32'h820FFFF2;
rContents[496] = 32'h41E00000;
rContents[497] = 32'h41D00000;
rContents[498] = 32'h41C00000;
rContents[499] = 32'hF0000000;
rContents[500] = 32'h61C00000;
rContents[501] = 32'h61D00000;
rContents[502] = 32'h61E00000;
rContents[503] = 32'h18111004;
rContents[504] = 32'h41D00000;
rContents[505] = 32'h41C00000;
rContents[506] = 32'h18011006;
rContents[507] = 32'h08ED0000;
rContents[508] = 32'h187DD002;
rContents[509] = 32'h100CCD00;
rContents[510] = 32'h4CF00000;
rContents[511] = 32'h2D000003;
rContents[512] = 32'h182EE003;
rContents[513] = 32'h101EDE00;
rContents[514] = 32'h186EE003;
rContents[515] = 32'h10DFFEFF;
rContents[516] = 32'h41E00000;
rContents[517] = 32'h41D00000;
rContents[518] = 32'h41C00000;
rContents[519] = 32'hF0000000;
rContents[520] = 32'h61C00000;
rContents[521] = 32'h61D00000;
rContents[522] = 32'h18111003;
rContents[523] = 32'h2D000000;
rContents[524] = 32'h41C00000;
rContents[525] = 32'h18011004;
rContents[526] = 32'h61C00000;
rContents[527] = 32'h61D00000;
rContents[528] = 32'hD00FFFE4;
rContents[529] = 32'h41D00000;
rContents[530] = 32'h18E0F000;
rContents[531] = 32'h81000007;
rContents[532] = 32'h61F00000;
rContents[533] = 32'hD00FFF29;
rContents[534] = 32'hD00001B5;
rContents[535] = 32'h41F00000;
rContents[536] = 32'h180DD001;
rContents[537] = 32'h800FFFF6;
rContents[538] = 32'h41C00000;
rContents[539] = 32'h41D00000;
rContents[540] = 32'h41C00000;
rContents[541] = 32'hF0000000;
rContents[542] = 32'h61C00000;
rContents[543] = 32'h61D00000;
rContents[544] = 32'h61E00000;
rContents[545] = 32'h2C000000;
rContents[546] = 32'h61C00000;
rContents[547] = 32'hD00FFF63;
rContents[548] = 32'h41C00000;
rContents[549] = 32'h2C00000B;
rContents[550] = 32'hD00FFF96;
rContents[551] = 32'h181CC001;
rContents[552] = 32'h18E0C000;
rContents[553] = 32'h820FFFFD;
rContents[554] = 32'h2C000001;
rContents[555] = 32'h61C00000;
rContents[556] = 32'hD00FFF5A;
rContents[557] = 32'h41C00000;
rContents[558] = 32'h2C000000;
rContents[559] = 32'h61C00000;
rContents[560] = 32'h2C000000;
rContents[561] = 32'h61C00000;
rContents[562] = 32'h2D000001;
rContents[563] = 32'h186DD000;
rContents[564] = 32'h2E000000;
rContents[565] = 32'hD0000084;
rContents[566] = 32'h10E0FD00;
rContents[567] = 32'h81000005;
rContents[568] = 32'h180EE001;
rContents[569] = 32'h18E0E402;
rContents[570] = 32'h8100006E;
rContents[571] = 32'h800FFFFA;
rContents[572] = 32'h41C00000;
rContents[573] = 32'h41C00000;
rContents[574] = 32'h2C000008;
rContents[575] = 32'h61C00000;
rContents[576] = 32'h2C0001AA;
rContents[577] = 32'h61C00000;
rContents[578] = 32'hD0000077;
rContents[579] = 32'h41C00000;
rContents[580] = 32'h41C00000;
rContents[581] = 32'h2D000001;
rContents[582] = 32'h186DD002;
rContents[583] = 32'h10F0FD00;
rContents[584] = 32'h8200000C;
rContents[585] = 32'hD00FFF73;
rContents[586] = 32'hD00FFF72;
rContents[587] = 32'hD00FFF71;
rContents[588] = 32'h18F0F001;
rContents[589] = 32'h8100005D;
rContents[590] = 32'hD00FFF6E;
rContents[591] = 32'h18E0F0AA;
rContents[592] = 32'h8200005A;
rContents[593] = 32'h2E000001;
rContents[594] = 32'h186EE001;
rContents[595] = 32'h80000014;
rContents[596] = 32'h2C000037;
rContents[597] = 32'h61C00000;
rContents[598] = 32'h2C000000;
rContents[599] = 32'h61C00000;
rContents[600] = 32'hD0000061;
rContents[601] = 32'h41C00000;
rContents[602] = 32'h41C00000;
rContents[603] = 32'h2C000029;
rContents[604] = 32'h61C00000;
rContents[605] = 32'h2C000000;
rContents[606] = 32'h61C00000;
rContents[607] = 32'hD000005A;
rContents[608] = 32'h41C00000;
rContents[609] = 32'h41C00000;
rContents[610] = 32'h2E000000;
rContents[611] = 32'h10E0FD00;
rContents[612] = 32'h82000003;
rContents[613] = 32'h2E000001;
rContents[614] = 32'h186EE000;
rContents[615] = 32'h2D000000;
rContents[616] = 32'h18F0E003;
rContents[617] = 32'h81000013;
rContents[618] = 32'h2C000037;
rContents[619] = 32'h61C00000;
rContents[620] = 32'h2C000000;
rContents[621] = 32'h61C00000;
rContents[622] = 32'hD000004B;
rContents[623] = 32'h41C00000;
rContents[624] = 32'h41C00000;
rContents[625] = 32'h2C000029;
rContents[626] = 32'h61C00000;
rContents[627] = 32'h2C000000;
rContents[628] = 32'h18F0E002;
rContents[629] = 32'h81000002;
rContents[630] = 32'h2C804000;
rContents[631] = 32'h61C00000;
rContents[632] = 32'hD0000041;
rContents[633] = 32'h41C00000;
rContents[634] = 32'h41C00000;
rContents[635] = 32'h80000008;
rContents[636] = 32'h2C000029;
rContents[637] = 32'h61C00000;
rContents[638] = 32'h2C000000;
rContents[639] = 32'h61C00000;
rContents[640] = 32'hD0000039;
rContents[641] = 32'h41C00000;
rContents[642] = 32'h41C00000;
rContents[643] = 32'h18F0F001;
rContents[644] = 32'h81000005;
rContents[645] = 32'h180DD001;
rContents[646] = 32'h18E0D480;
rContents[647] = 32'h81000023;
rContents[648] = 32'h800FFFE0;
rContents[649] = 32'h18F0E002;
rContents[650] = 32'h81000013;
rContents[651] = 32'h2C00003A;
rContents[652] = 32'h61C00000;
rContents[653] = 32'h2C000000;
rContents[654] = 32'h61C00000;
rContents[655] = 32'hD000002A;
rContents[656] = 32'h41C00000;
rContents[657] = 32'h41C00000;
rContents[658] = 32'h18E0F000;
rContents[659] = 32'h82000017;
rContents[660] = 32'hD00FFF28;
rContents[661] = 32'h18F0F040;
rContents[662] = 32'h81000004;
rContents[663] = 32'h2C000001;
rContents[664] = 32'h186CC002;
rContents[665] = 32'h103EEC00;
rContents[666] = 32'hD00FFF22;
rContents[667] = 32'hD00FFF21;
rContents[668] = 32'hD00FFF20;
rContents[669] = 32'h2C000010;
rContents[670] = 32'h61C00000;
rContents[671] = 32'h2C000200;
rContents[672] = 32'h61C00000;
rContents[673] = 32'hD0000018;
rContents[674] = 32'h41C00000;
rContents[675] = 32'h41C00000;
rContents[676] = 32'h18E0F000;
rContents[677] = 32'h82000005;
rContents[678] = 32'h8000000A;
rContents[679] = 32'hD00001AB;
rContents[680] = 32'h41C00000;
rContents[681] = 32'h41C00000;
rContents[682] = 32'h2C000000;
rContents[683] = 32'h61C00000;
rContents[684] = 32'hD00FFEDA;
rContents[685] = 32'h41C00000;
rContents[686] = 32'h2F0000FF;
rContents[687] = 32'h80000006;
rContents[688] = 32'h2C000000;
rContents[689] = 32'h61C00000;
rContents[690] = 32'hD00FFED4;
rContents[691] = 32'h41C00000;
rContents[692] = 32'h08FE0000;
rContents[693] = 32'h41E00000;
rContents[694] = 32'h41D00000;
rContents[695] = 32'h41C00000;
rContents[696] = 32'hF0000000;
rContents[697] = 32'h61C00000;
rContents[698] = 32'h61D00000;
rContents[699] = 32'h18111003;
rContents[700] = 32'h41D00000;
rContents[701] = 32'h41C00000;
rContents[702] = 32'h18011005;
rContents[703] = 32'hD00FFEFD;
rContents[704] = 32'h183CC040;
rContents[705] = 32'h61C00000;
rContents[706] = 32'hD00FFED8;
rContents[707] = 32'h41C00000;
rContents[708] = 32'h61C00000;
rContents[709] = 32'h08CD0000;
rContents[710] = 32'h18DDCCFF;
rContents[711] = 32'h61D00000;
rContents[712] = 32'hD00FFED2;
rContents[713] = 32'h41D00000;
rContents[714] = 32'h18DDC8FF;
rContents[715] = 32'h61D00000;
rContents[716] = 32'hD00FFECE;
rContents[717] = 32'h41D00000;
rContents[718] = 32'h18DDC4FF;
rContents[719] = 32'h61D00000;
rContents[720] = 32'hD00FFECA;
rContents[721] = 32'h41D00000;
rContents[722] = 32'h18DDC0FF;
rContents[723] = 32'h61D00000;
rContents[724] = 32'hD00FFEC6;
rContents[725] = 32'h41D00000;
rContents[726] = 32'h41C00000;
rContents[727] = 32'h18E0C040;
rContents[728] = 32'h82000003;
rContents[729] = 32'h2D000095;
rContents[730] = 32'h80000006;
rContents[731] = 32'h18E0C048;
rContents[732] = 32'h82000003;
rContents[733] = 32'h2D000087;
rContents[734] = 32'h80000002;
rContents[735] = 32'h2D0000FF;
rContents[736] = 32'h61D00000;
rContents[737] = 32'hD00FFEB9;
rContents[738] = 32'h41D00000;
rContents[739] = 32'h2D00000A;
rContents[740] = 32'hD00FFED8;
rContents[741] = 32'h18E0F0FF;
rContents[742] = 32'h82000005;
rContents[743] = 32'h181DD001;
rContents[744] = 32'h18E0D000;
rContents[745] = 32'h81000002;
rContents[746] = 32'h800FFFFA;
rContents[747] = 32'h41D00000;
rContents[748] = 32'h41C00000;
rContents[749] = 32'hF0000000;
rContents[750] = 32'h61C00000;
rContents[751] = 32'h61D00000;
rContents[752] = 32'h61E00000;
rContents[753] = 32'h18111004;
rContents[754] = 32'h41D00000;
rContents[755] = 32'h41C00000;
rContents[756] = 32'h18011006;
rContents[757] = 32'h2F000001;
rContents[758] = 32'h61F00000;
rContents[759] = 32'hD00FFE8F;
rContents[760] = 32'h41F00000;
rContents[761] = 32'h2F000011;
rContents[762] = 32'h61F00000;
rContents[763] = 32'h61D00000;
rContents[764] = 32'hD00FFFBD;
rContents[765] = 32'h18111002;
rContents[766] = 32'h18E0F000;
rContents[767] = 32'h8200001E;
rContents[768] = 32'hD00FFEBC;
rContents[769] = 32'h18E0F0FE;
rContents[770] = 32'h820FFFFE;
rContents[771] = 32'h2E000080;
rContents[772] = 32'h2D000000;
rContents[773] = 32'hD00FFEB7;
rContents[774] = 32'h186DF018;
rContents[775] = 32'hD00FFEB5;
rContents[776] = 32'h186FF010;
rContents[777] = 32'h103DDF00;
rContents[778] = 32'hD00FFEB2;
rContents[779] = 32'h186FF008;
rContents[780] = 32'h103DDF00;
rContents[781] = 32'hD00FFEAF;
rContents[782] = 32'h103DDF00;
rContents[783] = 32'h6CD00000;
rContents[784] = 32'h180CC001;
rContents[785] = 32'h181EE001;
rContents[786] = 32'h18E0E000;
rContents[787] = 32'h820FFFF2;
rContents[788] = 32'hD00FFEA8;
rContents[789] = 32'hD00FFEA7;
rContents[790] = 32'h2F000000;
rContents[791] = 32'h61F00000;
rContents[792] = 32'hD00FFE6E;
rContents[793] = 32'h41F00000;
rContents[794] = 32'hD00FFEA2;
rContents[795] = 32'h2F000000;
rContents[796] = 32'h80000006;
rContents[797] = 32'h2F000000;
rContents[798] = 32'h61F00000;
rContents[799] = 32'hD00FFE67;
rContents[800] = 32'h41F00000;
rContents[801] = 32'h2F0000FF;
rContents[802] = 32'h41E00000;
rContents[803] = 32'h41D00000;
rContents[804] = 32'h41C00000;
rContents[805] = 32'hF0000000;
rContents[806] = 32'h61C00000;
rContents[807] = 32'h61D00000;
rContents[808] = 32'h61E00000;
rContents[809] = 32'h18111004;
rContents[810] = 32'h41D00000;
rContents[811] = 32'h41C00000;
rContents[812] = 32'h18011006;
rContents[813] = 32'h2F000001;
rContents[814] = 32'h61F00000;
rContents[815] = 32'hD00FFE57;
rContents[816] = 32'h41F00000;
rContents[817] = 32'h2F000018;
rContents[818] = 32'h61F00000;
rContents[819] = 32'h61D00000;
rContents[820] = 32'hD00FFF85;
rContents[821] = 32'h18111002;
rContents[822] = 32'h18E0F000;
rContents[823] = 32'h8200002E;
rContents[824] = 32'h2F0000FE;
rContents[825] = 32'h61F00000;
rContents[826] = 32'hD00FFE60;
rContents[827] = 32'h41F00000;
rContents[828] = 32'h2E000080;
rContents[829] = 32'h4CD00000;
rContents[830] = 32'h61C00000;
rContents[831] = 32'h182CDCFF;
rContents[832] = 32'h188DD018;
rContents[833] = 32'h61D00000;
rContents[834] = 32'hD00FFE58;
rContents[835] = 32'h41D00000;
rContents[836] = 32'h182CD8FF;
rContents[837] = 32'h188DD010;
rContents[838] = 32'h61D00000;
rContents[839] = 32'hD00FFE53;
rContents[840] = 32'h41D00000;
rContents[841] = 32'h182CD4FF;
rContents[842] = 32'h188DD008;
rContents[843] = 32'h61D00000;
rContents[844] = 32'hD00FFE4E;
rContents[845] = 32'h41D00000;
rContents[846] = 32'h182CD0FF;
rContents[847] = 32'h61D00000;
rContents[848] = 32'hD00FFE4A;
rContents[849] = 32'h41D00000;
rContents[850] = 32'h41C00000;
rContents[851] = 32'h180CC001;
rContents[852] = 32'h181EE001;
rContents[853] = 32'h18E0E000;
rContents[854] = 32'h820FFFE7;
rContents[855] = 32'h2F0000FF;
rContents[856] = 32'h61F00000;
rContents[857] = 32'hD00FFE41;
rContents[858] = 32'hD00FFE40;
rContents[859] = 32'h41F00000;
rContents[860] = 32'hD00FFE60;
rContents[861] = 32'h18E0F0FF;
rContents[862] = 32'h820FFFFE;
rContents[863] = 32'h2F000000;
rContents[864] = 32'h61F00000;
rContents[865] = 32'hD00FFE25;
rContents[866] = 32'h41F00000;
rContents[867] = 32'h2F000000;
rContents[868] = 32'h80000006;
rContents[869] = 32'h2F000000;
rContents[870] = 32'h61F00000;
rContents[871] = 32'hD00FFE1F;
rContents[872] = 32'h41F00000;
rContents[873] = 32'h2F0000FF;
rContents[874] = 32'h41E00000;
rContents[875] = 32'h41D00000;
rContents[876] = 32'h41C00000;
rContents[877] = 32'hF0000000;
rContents[878] = 32'h61D00000;
rContents[879] = 32'h2D000030;
rContents[880] = 32'h61D00000;
rContents[881] = 32'h2D000000;
rContents[882] = 32'h61D00000;
rContents[883] = 32'hD00FFD98;
rContents[884] = 32'h41D00000;
rContents[885] = 32'h41D00000;
rContents[886] = 32'h2D000031;
rContents[887] = 32'h61D00000;
rContents[888] = 32'h2D000000;
rContents[889] = 32'h61D00000;
rContents[890] = 32'hD00FFD91;
rContents[891] = 32'h41D00000;
rContents[892] = 32'h41D00000;
rContents[893] = 32'h2D000032;
rContents[894] = 32'h61D00000;
rContents[895] = 32'h2D000000;
rContents[896] = 32'h61D00000;
rContents[897] = 32'hD00FFD8A;
rContents[898] = 32'h41D00000;
rContents[899] = 32'h41D00000;
rContents[900] = 32'hD0000003;
rContents[901] = 32'h41D00000;
rContents[902] = 32'hF0000000;
rContents[903] = 32'h61D00000;
rContents[904] = 32'h2D000031;
rContents[905] = 32'h61D00000;
rContents[906] = 32'h2D000000;
rContents[907] = 32'h61D00000;
rContents[908] = 32'hD00FFD7F;
rContents[909] = 32'h41D00000;
rContents[910] = 32'h41D00000;
rContents[911] = 32'h2D000032;
rContents[912] = 32'h61D00000;
rContents[913] = 32'h2D000000;
rContents[914] = 32'h61D00000;
rContents[915] = 32'hD00FFD78;
rContents[916] = 32'h41D00000;
rContents[917] = 32'h41D00000;
rContents[918] = 32'h2D000033;
rContents[919] = 32'h61D00000;
rContents[920] = 32'h2D000000;
rContents[921] = 32'h61D00000;
rContents[922] = 32'hD00FFD71;
rContents[923] = 32'h41D00000;
rContents[924] = 32'h41D00000;
rContents[925] = 32'h2D000031;
rContents[926] = 32'h61D00000;
rContents[927] = 32'hD00FFD83;
rContents[928] = 32'h41D00000;
rContents[929] = 32'h180FF001;
rContents[930] = 32'h61F00000;
rContents[931] = 32'h2D000031;
rContents[932] = 32'h61D00000;
rContents[933] = 32'h61F00000;
rContents[934] = 32'hD00FFD65;
rContents[935] = 32'h41F00000;
rContents[936] = 32'h41D00000;
rContents[937] = 32'h41F00000;
rContents[938] = 32'h18E0F050;
rContents[939] = 32'h820FFFEB;
rContents[940] = 32'h2D000031;
rContents[941] = 32'h61D00000;
rContents[942] = 32'h2D000000;
rContents[943] = 32'h61D00000;
rContents[944] = 32'hD00FFD5B;
rContents[945] = 32'h41D00000;
rContents[946] = 32'h41D00000;
rContents[947] = 32'h2D000032;
rContents[948] = 32'h61D00000;
rContents[949] = 32'hD00FFD6D;
rContents[950] = 32'h41D00000;
rContents[951] = 32'h180FF001;
rContents[952] = 32'h61F00000;
rContents[953] = 32'h2D000032;
rContents[954] = 32'h61D00000;
rContents[955] = 32'h61F00000;
rContents[956] = 32'hD00FFD4F;
rContents[957] = 32'h41F00000;
rContents[958] = 32'h41D00000;
rContents[959] = 32'h41F00000;
rContents[960] = 32'h18E0F028;
rContents[961] = 32'h820FFFD5;
rContents[962] = 32'h2D000032;
rContents[963] = 32'h61D00000;
rContents[964] = 32'h2D000000;
rContents[965] = 32'h61D00000;
rContents[966] = 32'hD00FFD45;
rContents[967] = 32'h41D00000;
rContents[968] = 32'h41D00000;
rContents[969] = 32'h41D00000;
rContents[970] = 32'hF0000000;
rContents[971] = 32'h61C00000;
rContents[972] = 32'h61D00000;
rContents[973] = 32'h18111003;
rContents[974] = 32'h41C00000;
rContents[975] = 32'h18011004;
rContents[976] = 32'h18E0C020;
rContents[977] = 32'h8300001E;
rContents[978] = 32'h18E0C00D;
rContents[979] = 32'h82000009;
rContents[980] = 32'h2D000031;
rContents[981] = 32'h61D00000;
rContents[982] = 32'h2D000000;
rContents[983] = 32'h61D00000;
rContents[984] = 32'hD00FFD33;
rContents[985] = 32'h41D00000;
rContents[986] = 32'h41D00000;
rContents[987] = 32'h80000048;
rContents[988] = 32'h18E0C00A;
rContents[989] = 32'h82000011;
rContents[990] = 32'h2D000032;
rContents[991] = 32'h61D00000;
rContents[992] = 32'hD00FFD42;
rContents[993] = 32'h41D00000;
rContents[994] = 32'h180FF001;
rContents[995] = 32'h61F00000;
rContents[996] = 32'h2D000032;
rContents[997] = 32'h61D00000;
rContents[998] = 32'h61F00000;
rContents[999] = 32'hD00FFD24;
rContents[1000] = 32'h41F00000;
rContents[1001] = 32'h41D00000;
rContents[1002] = 32'h41F00000;
rContents[1003] = 32'h18E0F028;
rContents[1004] = 32'h81000036;
rContents[1005] = 32'h80000036;
rContents[1006] = 32'h80000035;
rContents[1007] = 32'h183CC4FF;
rContents[1008] = 32'h2D000033;
rContents[1009] = 32'h61D00000;
rContents[1010] = 32'h61C00000;
rContents[1011] = 32'hD00FFD18;
rContents[1012] = 32'h41C00000;
rContents[1013] = 32'h41D00000;
rContents[1014] = 32'h2D000031;
rContents[1015] = 32'h61D00000;
rContents[1016] = 32'hD00FFD2A;
rContents[1017] = 32'h41D00000;
rContents[1018] = 32'h180FF001;
rContents[1019] = 32'h61F00000;
rContents[1020] = 32'h2D000031;
rContents[1021] = 32'h61D00000;
rContents[1022] = 32'h61F00000;
rContents[1023] = 32'hD00FFD0C;
rContents[1024] = 32'h41F00000;
rContents[1025] = 32'h41D00000;
rContents[1026] = 32'h41F00000;
rContents[1027] = 32'h18E0F050;
rContents[1028] = 32'h8200001F;
rContents[1029] = 32'h2D000031;
rContents[1030] = 32'h61D00000;
rContents[1031] = 32'h2D000000;
rContents[1032] = 32'h61D00000;
rContents[1033] = 32'hD00FFD02;
rContents[1034] = 32'h41D00000;
rContents[1035] = 32'h41D00000;
rContents[1036] = 32'h2D000032;
rContents[1037] = 32'h61D00000;
rContents[1038] = 32'hD00FFD14;
rContents[1039] = 32'h41D00000;
rContents[1040] = 32'h180FF001;
rContents[1041] = 32'h61F00000;
rContents[1042] = 32'h2D000032;
rContents[1043] = 32'h61D00000;
rContents[1044] = 32'h61F00000;
rContents[1045] = 32'hD00FFCF6;
rContents[1046] = 32'h41F00000;
rContents[1047] = 32'h41D00000;
rContents[1048] = 32'h41F00000;
rContents[1049] = 32'h18E0F028;
rContents[1050] = 32'h82000009;
rContents[1051] = 32'h2D000032;
rContents[1052] = 32'h61D00000;
rContents[1053] = 32'h2D000000;
rContents[1054] = 32'h61D00000;
rContents[1055] = 32'hD00FFCEC;
rContents[1056] = 32'h41D00000;
rContents[1057] = 32'h41D00000;
rContents[1058] = 32'hD00FFF65;
rContents[1059] = 32'h41D00000;
rContents[1060] = 32'h41C00000;
rContents[1061] = 32'hF0000000;
rContents[1062] = 32'h0A0A416E;
rContents[1063] = 32'h20657272;
rContents[1064] = 32'h6F722068;
rContents[1065] = 32'h6173206F;
rContents[1066] = 32'h63637572;
rContents[1067] = 32'h65642E0A;
rContents[1068] = 32'h00000000;
rContents[1069] = 32'h0A0A4120;
rContents[1070] = 32'h66617461;
rContents[1071] = 32'h6C206572;
rContents[1072] = 32'h726F7220;
rContents[1073] = 32'h68617320;
rContents[1074] = 32'h6F636375;
rContents[1075] = 32'h7265642E;
rContents[1076] = 32'h0A000000;
rContents[1077] = 32'h43616C6C;
rContents[1078] = 32'h65642061;
rContents[1079] = 32'h74200000;
rContents[1080] = 32'h53746163;
rContents[1081] = 32'h6B747261;
rContents[1082] = 32'h63652028;
rContents[1083] = 32'h746F7020;
rContents[1084] = 32'h3136293A;
rContents[1085] = 32'h0A000000;
rContents[1086] = 32'h52656769;
rContents[1087] = 32'h73746572;
rContents[1088] = 32'h733A0A00;
rContents[1089] = 32'h52657375;
rContents[1090] = 32'h6D696E67;
rContents[1091] = 32'h2E0A0A00;
rContents[1092] = 32'h48616C74;
rContents[1093] = 32'h696E672E;
rContents[1094] = 32'h0A0A0000;
rContents[1095] = 32'h80000001;
rContents[1096] = 32'h2F00042D;
rContents[1097] = 32'h61F00000;
rContents[1098] = 32'hD00FFDBE;
rContents[1099] = 32'h41F00000;
rContents[1100] = 32'h2F000435;
rContents[1101] = 32'h61F00000;
rContents[1102] = 32'hD00FFDBA;
rContents[1103] = 32'h41F00000;
rContents[1104] = 32'hD00FFD8A;
rContents[1105] = 32'h04200000;
rContents[1106] = 32'h61F00000;
rContents[1107] = 32'h2F000435;
rContents[1108] = 32'h61F00000;
rContents[1109] = 32'hD00FFDB3;
rContents[1110] = 32'h41F00000;
rContents[1111] = 32'h2F0000F0;
rContents[1112] = 32'h181FF001;
rContents[1113] = 32'h18E0F000;
rContents[1114] = 32'h820FFFFE;
rContents[1115] = 32'h18111001;
rContents[1116] = 32'hD00FFD7E;
rContents[1117] = 32'h18011001;
rContents[1118] = 32'h2F00000A;
rContents[1119] = 32'h61F00000;
rContents[1120] = 32'hD0000013;
rContents[1121] = 32'h41F00000;
rContents[1122] = 32'h2F00000D;
rContents[1123] = 32'h61F00000;
rContents[1124] = 32'hD000000F;
rContents[1125] = 32'h41F00000;
rContents[1126] = 32'h41F00000;
rContents[1127] = 32'hF0000000;
rContents[1128] = 32'hF0000000;
rContents[1129] = 32'hF0000000;
rContents[1130] = 32'h4C656D6F;
rContents[1131] = 32'h6E207630;
rContents[1132] = 32'h2E32202D;
rContents[1133] = 32'h20666F72;
rContents[1134] = 32'h20657052;
rContents[1135] = 32'h49534320;
rContents[1136] = 32'h76352073;
rContents[1137] = 32'h79737465;
rContents[1138] = 32'h6D730000;
rContents[1139] = 32'h18111001;
rContents[1140] = 32'h41F00000;
rContents[1141] = 32'h18011002;
rContents[1142] = 32'h61F00000;
rContents[1143] = 32'hD00FFCC7;
rContents[1144] = 32'hD00FFF53;
rContents[1145] = 32'h41F00000;
rContents[1146] = 32'hF0000000;
rContents[1147] = 32'h800FFCDF;
rContents[1148] = 32'h800FFD5E;
rContents[1149] = 32'h800FFD8B;
rContents[1150] = 32'h800FFFCA;
rContents[1151] = 32'h210017FF;
rContents[1152] = 32'h2800046A;
rContents[1153] = 32'h61800000;
rContents[1154] = 32'hD00FFFFB;
rContents[1155] = 32'h41800000;
rContents[1156] = 32'h26001000;
rContents[1157] = 32'h29000000;
rContents[1158] = 32'h2800000A;
rContents[1159] = 32'h61800000;
rContents[1160] = 32'hD00FFFEB;
rContents[1161] = 32'h41800000;
rContents[1162] = 32'h2800000D;
rContents[1163] = 32'h61800000;
rContents[1164] = 32'hD00FFFE7;
rContents[1165] = 32'h41800000;
rContents[1166] = 32'h2800003E;
rContents[1167] = 32'h61800000;
rContents[1168] = 32'hD00FFFE3;
rContents[1169] = 32'h41800000;
rContents[1170] = 32'hD00FFFE9;
rContents[1171] = 32'h18E0F008;
rContents[1172] = 32'h8200000E;
rContents[1173] = 32'h18E06000;
rContents[1174] = 32'h82000002;
rContents[1175] = 32'h800FFFFB;
rContents[1176] = 32'h18166002;
rContents[1177] = 32'h18199001;
rContents[1178] = 32'h46F00000;
rContents[1179] = 32'h61F00000;
rContents[1180] = 32'hD00FFFD7;
rContents[1181] = 32'h41F00000;
rContents[1182] = 32'h18066001;
rContents[1183] = 32'h2F000000;
rContents[1184] = 32'h66F00000;
rContents[1185] = 32'h800FFFF1;
rContents[1186] = 32'h18E0F00D;
rContents[1187] = 32'h82000003;
rContents[1188] = 32'h66F00000;
rContents[1189] = 32'h8000000A;
rContents[1190] = 32'h18F09180;
rContents[1191] = 32'h820FFFEB;
rContents[1192] = 32'h61F00000;
rContents[1193] = 32'hD00FFFCA;
rContents[1194] = 32'h41F00000;
rContents[1195] = 32'h66F00000;
rContents[1196] = 32'h18066001;
rContents[1197] = 32'h18099001;
rContents[1198] = 32'h800FFFE4;
rContents[1199] = 32'h26001000;
rContents[1200] = 32'h27000000;
rContents[1201] = 32'h46900000;
rContents[1202] = 32'h18E0900D;
rContents[1203] = 32'h82000005;
rContents[1204] = 32'h18E0703A;
rContents[1205] = 32'h82000002;
rContents[1206] = 32'h41800000;
rContents[1207] = 32'h800FFFCD;
rContents[1208] = 32'h18E09052;
rContents[1209] = 32'h8200000C;
rContents[1210] = 32'h2800000A;
rContents[1211] = 32'h61800000;
rContents[1212] = 32'hD00FFFB7;
rContents[1213] = 32'h41800000;
rContents[1214] = 32'h2800000D;
rContents[1215] = 32'h61800000;
rContents[1216] = 32'hD00FFFB3;
rContents[1217] = 32'h41800000;
rContents[1218] = 32'hD0400000;
rContents[1219] = 32'h18066001;
rContents[1220] = 32'h800FFFED;
rContents[1221] = 32'h18E0903A;
rContents[1222] = 32'h82000005;
rContents[1223] = 32'h2700003A;
rContents[1224] = 32'h61400000;
rContents[1225] = 32'h18066001;
rContents[1226] = 32'h800FFFE7;
rContents[1227] = 32'h18E0902E;
rContents[1228] = 32'h82000007;
rContents[1229] = 32'h18E0703A;
rContents[1230] = 32'h82000002;
rContents[1231] = 32'h41800000;
rContents[1232] = 32'h2700002E;
rContents[1233] = 32'h18066001;
rContents[1234] = 32'h800FFFDF;
rContents[1235] = 32'h18E09020;
rContents[1236] = 32'h82000003;
rContents[1237] = 32'h18066001;
rContents[1238] = 32'h800FFFDB;
rContents[1239] = 32'h25000000;
rContents[1240] = 32'h46900000;
rContents[1241] = 32'h18199030;
rContents[1242] = 32'h18E0900A;
rContents[1243] = 32'h84000007;
rContents[1244] = 32'h18199007;
rContents[1245] = 32'h18E0900A;
rContents[1246] = 32'h84000008;
rContents[1247] = 32'h18E09010;
rContents[1248] = 32'h84000002;
rContents[1249] = 32'h80000005;
rContents[1250] = 32'h18655004;
rContents[1251] = 32'h10355900;
rContents[1252] = 32'h18066001;
rContents[1253] = 32'h800FFFF3;
rContents[1254] = 32'h46900000;
rContents[1255] = 32'h18E0703A;
rContents[1256] = 32'h82000004;
rContents[1257] = 32'h64500000;
rContents[1258] = 32'h18044001;
rContents[1259] = 32'h800FFFC6;
rContents[1260] = 32'h61400000;
rContents[1261] = 32'h08450000;
rContents[1262] = 32'h18E0902E;
rContents[1263] = 32'h82000003;
rContents[1264] = 32'h41800000;
rContents[1265] = 32'h800FFFC0;
rContents[1266] = 32'h18E07000;
rContents[1267] = 32'h82000016;
rContents[1268] = 32'h41800000;
rContents[1269] = 32'h2800000A;
rContents[1270] = 32'h61800000;
rContents[1271] = 32'hD00FFF7C;
rContents[1272] = 32'h41800000;
rContents[1273] = 32'h2800000D;
rContents[1274] = 32'h61800000;
rContents[1275] = 32'hD00FFF78;
rContents[1276] = 32'h41800000;
rContents[1277] = 32'h61400000;
rContents[1278] = 32'hD00FFCDC;
rContents[1279] = 32'h41400000;
rContents[1280] = 32'h2800003A;
rContents[1281] = 32'h61800000;
rContents[1282] = 32'hD00FFF71;
rContents[1283] = 32'h41800000;
rContents[1284] = 32'h44800000;
rContents[1285] = 32'h61800000;
rContents[1286] = 32'hD00FFF76;
rContents[1287] = 32'h41800000;
rContents[1288] = 32'h800FFFA9;
rContents[1289] = 32'h18E0702E;
rContents[1290] = 32'hD20FFF74;
rContents[1291] = 32'h08840000;
rContents[1292] = 32'h41400000;
rContents[1293] = 32'h10E08400;
rContents[1294] = 32'h8B000002;
rContents[1295] = 32'h08840000;
rContents[1296] = 32'h101A8400;
rContents[1297] = 32'h180AA001;
rContents[1298] = 32'h61400000;
rContents[1299] = 32'h2800000A;
rContents[1300] = 32'h61800000;
rContents[1301] = 32'hD00FFF5E;
rContents[1302] = 32'h41800000;
rContents[1303] = 32'h2800000D;
rContents[1304] = 32'h61800000;
rContents[1305] = 32'hD00FFF5A;
rContents[1306] = 32'h41800000;
rContents[1307] = 32'h61400000;
rContents[1308] = 32'hD00FFCBE;
rContents[1309] = 32'h41400000;
rContents[1310] = 32'h2800003A;
rContents[1311] = 32'h61800000;
rContents[1312] = 32'hD00FFF53;
rContents[1313] = 32'h41800000;
rContents[1314] = 32'h18E0A008;
rContents[1315] = 32'h83000003;
rContents[1316] = 32'h08BA0000;
rContents[1317] = 32'h80000002;
rContents[1318] = 32'h2B000008;
rContents[1319] = 32'h101AAB00;
rContents[1320] = 32'h28000020;
rContents[1321] = 32'h61800000;
rContents[1322] = 32'hD00FFF49;
rContents[1323] = 32'h41800000;
rContents[1324] = 32'h44800000;
rContents[1325] = 32'h61800000;
rContents[1326] = 32'hD00FFF4E;
rContents[1327] = 32'h41800000;
rContents[1328] = 32'h18044001;
rContents[1329] = 32'h181BB001;
rContents[1330] = 32'h18E0B000;
rContents[1331] = 32'h820FFFF5;
rContents[1332] = 32'h18E0A000;
rContents[1333] = 32'h820FFFDE;
rContents[1334] = 32'h41400000;
rContents[1335] = 32'h27000000;
rContents[1336] = 32'h800FFF79;
    end

endmodule

/*  Program 1 - square wave generator over GPIO
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808000;
        rContents[8] = 32'h3500FFFF;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25000000;
        rContents[17] = 32'h08650000;
        rContents[18] = 32'h36808002;
        rContents[19] = 32'h64600001;
        rContents[20] = 32'h27010005;
        rContents[21] = 32'h64700000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h04000000;
        rContents[26] = 32'h18B5580F;
        rContents[27] = 32'h18055001;
        rContents[28] = 32'h800FFFF5;
        rContents[29] = 32'h0;
        rContents[30] = 32'h0;
        rContents[31] = 32'h0;
        rContents[32] = 32'h0;
        rContents[33] = 32'h0;
        rContents[34] = 32'h0;
        rContents[35] = 32'h0; */
        
/*  Program 2 - print some 'H's over the serial link
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808101;
        rContents[8] = 32'h35000048;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25808100;
        rContents[17] = 32'h35000080;
        rContents[18] = 32'h64500001;
        rContents[19] = 32'h27010005;
        rContents[20] = 32'h64700000;
        rContents[21] = 32'h04000000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h800FFFED; */
