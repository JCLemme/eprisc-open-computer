module epRISC_embeddedROM(iClk, iAddr, oData, iEnable);

    input iClk, iEnable;
    input [9:0] iAddr;
    output wire [31:0] oData;
    
    reg [31:0] rDataOut, rContents[0:1023];
    
    assign oData = (iEnable) ? rDataOut : 32'bz;
    
    always @(posedge iClk) begin
        rDataOut = rContents[iAddr];
    end
    
    initial begin
rContents[0] = 32'h21000410;
rContents[1] = 32'hD0000027;
rContents[2] = 32'h240034EA;
rContents[3] = 32'h24000201;
rContents[4] = 32'h61400000;
rContents[5] = 32'h24000000;
rContents[6] = 32'h61400000;
rContents[7] = 32'hD000002B;
rContents[8] = 32'h41400000;
rContents[9] = 32'h41400000;
rContents[10] = 32'h24000200;
rContents[11] = 32'h61400000;
rContents[12] = 32'h24000080;
rContents[13] = 32'h61400000;
rContents[14] = 32'hD0000024;
rContents[15] = 32'h41400000;
rContents[16] = 32'h41400000;
rContents[17] = 32'h04200000;
rContents[18] = 32'hD000007D;
rContents[19] = 32'h61F00000;
rContents[20] = 32'hD0000051;
rContents[21] = 32'h2400003A;
rContents[22] = 32'h61400000;
rContents[23] = 32'hD000004E;
rContents[24] = 32'h41400000;
rContents[25] = 32'h24000020;
rContents[26] = 32'h61400000;
rContents[27] = 32'hD000004A;
rContents[28] = 32'h41400000;
rContents[29] = 32'hD000009E;
rContents[30] = 32'h41F00000;
rContents[31] = 32'h2500000A;
rContents[32] = 32'h61500000;
rContents[33] = 32'hD0000044;
rContents[34] = 32'h41F00000;
rContents[35] = 32'h2500000D;
rContents[36] = 32'h61500000;
rContents[37] = 32'hD0000040;
rContents[38] = 32'h41F00000;
rContents[39] = 32'h800FFFEB;
rContents[40] = 32'h61C00000;
rContents[41] = 32'h2C000800;
rContents[42] = 32'h2F010001;
rContents[43] = 32'h6CF00000;
rContents[44] = 32'h04000000;
rContents[45] = 32'h04000000;
rContents[46] = 32'h04000000;
rContents[47] = 32'h04000000;
rContents[48] = 32'h41C00000;
rContents[49] = 32'hF0000000;
rContents[50] = 32'h61E00000;
rContents[51] = 32'h61D00000;
rContents[52] = 32'h61C00000;
rContents[53] = 32'h18111004;
rContents[54] = 32'h2C000800;
rContents[55] = 32'h41D00000;
rContents[56] = 32'h41E00000;
rContents[57] = 32'h2F600008;
rContents[58] = 32'h103FFE00;
rContents[59] = 32'h186FF010;
rContents[60] = 32'h103FFD00;
rContents[61] = 32'h6CF00001;
rContents[62] = 32'h2F010005;
rContents[63] = 32'h6CF00000;
rContents[64] = 32'h4CF00000;
rContents[65] = 32'h18F0F001;
rContents[66] = 32'h820FFFFE;
rContents[67] = 32'h4CF00002;
rContents[68] = 32'h18011006;
rContents[69] = 32'h41C00000;
rContents[70] = 32'h41D00000;
rContents[71] = 32'h41E00000;
rContents[72] = 32'hF0000000;
rContents[73] = 32'h61E00000;
rContents[74] = 32'h61C00000;
rContents[75] = 32'h18111003;
rContents[76] = 32'h2C000800;
rContents[77] = 32'h41E00000;
rContents[78] = 32'h2F600000;
rContents[79] = 32'h103FFE00;
rContents[80] = 32'h186FF010;
rContents[81] = 32'h6CF00001;
rContents[82] = 32'h2F010005;
rContents[83] = 32'h6CF00000;
rContents[84] = 32'h4CF00000;
rContents[85] = 32'h18F0F001;
rContents[86] = 32'h820FFFFE;
rContents[87] = 32'h2F600000;
rContents[88] = 32'h103FFE00;
rContents[89] = 32'h186FF010;
rContents[90] = 32'h6CF00001;
rContents[91] = 32'h2F010005;
rContents[92] = 32'h6CF00000;
rContents[93] = 32'h4CF00000;
rContents[94] = 32'h18F0F001;
rContents[95] = 32'h820FFFFE;
rContents[96] = 32'h4CF00002;
rContents[97] = 32'h18011004;
rContents[98] = 32'h41C00000;
rContents[99] = 32'h41E00000;
rContents[100] = 32'hF0000000;
rContents[101] = 32'h61D00000;
rContents[102] = 32'h61C00000;
rContents[103] = 32'h18111003;
rContents[104] = 32'h2C000800;
rContents[105] = 32'h41D00000;
rContents[106] = 32'h2F800100;
rContents[107] = 32'h6CF00001;
rContents[108] = 32'h2F010005;
rContents[109] = 32'h6CF00000;
rContents[110] = 32'h4CF00000;
rContents[111] = 32'h18F0F001;
rContents[112] = 32'h820FFFFE;
rContents[113] = 32'h2F800100;
rContents[114] = 32'h6CF00001;
rContents[115] = 32'h2F010005;
rContents[116] = 32'h6CF00000;
rContents[117] = 32'h4CF00000;
rContents[118] = 32'h18F0F001;
rContents[119] = 32'h820FFFFE;
rContents[120] = 32'h4CF00002;
rContents[121] = 32'h18F0F080;
rContents[122] = 32'h820FFFF7;
rContents[123] = 32'h2F808101;
rContents[124] = 32'h103FFD00;
rContents[125] = 32'h6CF00001;
rContents[126] = 32'h2F010005;
rContents[127] = 32'h6CF00000;
rContents[128] = 32'h4CF00000;
rContents[129] = 32'h18F0F001;
rContents[130] = 32'h820FFFFE;
rContents[131] = 32'h2F808100;
rContents[132] = 32'h3F000080;
rContents[133] = 32'h6CF00001;
rContents[134] = 32'h2F010005;
rContents[135] = 32'h6CF00000;
rContents[136] = 32'h4CF00000;
rContents[137] = 32'h18F0F001;
rContents[138] = 32'h820FFFFE;
rContents[139] = 32'h18011004;
rContents[140] = 32'h41C00000;
rContents[141] = 32'h41D00000;
rContents[142] = 32'hF0000000;
rContents[143] = 32'h61C00000;
rContents[144] = 32'h2C000800;
rContents[145] = 32'h2F808100;
rContents[146] = 32'h3F000020;
rContents[147] = 32'h6CF00001;
rContents[148] = 32'h2F010005;
rContents[149] = 32'h6CF00000;
rContents[150] = 32'h4CF00000;
rContents[151] = 32'h18F0F001;
rContents[152] = 32'h820FFFFE;
rContents[153] = 32'h2F800100;
rContents[154] = 32'h6CF00001;
rContents[155] = 32'h2F010005;
rContents[156] = 32'h6CF00000;
rContents[157] = 32'h4CF00000;
rContents[158] = 32'h18F0F001;
rContents[159] = 32'h820FFFFE;
rContents[160] = 32'h2F800100;
rContents[161] = 32'h6CF00001;
rContents[162] = 32'h2F010005;
rContents[163] = 32'h6CF00000;
rContents[164] = 32'h4CF00000;
rContents[165] = 32'h18F0F001;
rContents[166] = 32'h820FFFFE;
rContents[167] = 32'h4CF00002;
rContents[168] = 32'h18F0F020;
rContents[169] = 32'h820FFFF7;
rContents[170] = 32'h2F800102;
rContents[171] = 32'h6CF00001;
rContents[172] = 32'h2F010005;
rContents[173] = 32'h6CF00000;
rContents[174] = 32'h4CF00000;
rContents[175] = 32'h18F0F001;
rContents[176] = 32'h820FFFFE;
rContents[177] = 32'h2F800102;
rContents[178] = 32'h6CF00001;
rContents[179] = 32'h2F010005;
rContents[180] = 32'h6CF00000;
rContents[181] = 32'h4CF00000;
rContents[182] = 32'h18F0F001;
rContents[183] = 32'h820FFFFE;
rContents[184] = 32'h4CF00002;
rContents[185] = 32'h41C00000;
rContents[186] = 32'hF0000000;
rContents[187] = 32'h61C00000;
rContents[188] = 32'h61D00000;
rContents[189] = 32'h61E00000;
rContents[190] = 32'h18111004;
rContents[191] = 32'h41C00000;
rContents[192] = 32'h2E000008;
rContents[193] = 32'h18011005;
rContents[194] = 32'h182DCCF0;
rContents[195] = 32'h186CC004;
rContents[196] = 32'h188DD01C;
rContents[197] = 32'h180DD030;
rContents[198] = 32'h18E0D03A;
rContents[199] = 32'h83000002;
rContents[200] = 32'h180DD007;
rContents[201] = 32'h61D00000;
rContents[202] = 32'hD00FFF9B;
rContents[203] = 32'h41D00000;
rContents[204] = 32'h181EE001;
rContents[205] = 32'h18E0E000;
rContents[206] = 32'h8D0FFFF4;
rContents[207] = 32'h41E00000;
rContents[208] = 32'h41D00000;
rContents[209] = 32'h41C00000;
rContents[210] = 32'hF0000000;
    end

endmodule

/*  Program 1 - square wave generator over GPIO
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808000;
        rContents[8] = 32'h3500FFFF;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25000000;
        rContents[17] = 32'h08650000;
        rContents[18] = 32'h36808002;
        rContents[19] = 32'h64600001;
        rContents[20] = 32'h27010005;
        rContents[21] = 32'h64700000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h04000000;
        rContents[26] = 32'h18B5580F;
        rContents[27] = 32'h18055001;
        rContents[28] = 32'h800FFFF5;
        rContents[29] = 32'h0;
        rContents[30] = 32'h0;
        rContents[31] = 32'h0;
        rContents[32] = 32'h0;
        rContents[33] = 32'h0;
        rContents[34] = 32'h0;
        rContents[35] = 32'h0; */
        
/*  Program 2 - print some 'H's over the serial link
        rContents[0] = 32'h24000200;
        rContents[1] = 32'h27010001;
        rContents[2] = 32'h64700000;
        rContents[3] = 32'h04000000;
        rContents[4] = 32'h04000000;
        rContents[5] = 32'h04000000;
        rContents[6] = 32'h04000000;
        rContents[7] = 32'h25808101;
        rContents[8] = 32'h35000048;
        rContents[9] = 32'h64500001;
        rContents[10] = 32'h27010005;
        rContents[11] = 32'h64700000;
        rContents[12] = 32'h04000000;
        rContents[13] = 32'h04000000;
        rContents[14] = 32'h04000000;
        rContents[15] = 32'h04000000;
        rContents[16] = 32'h25808100;
        rContents[17] = 32'h35000080;
        rContents[18] = 32'h64500001;
        rContents[19] = 32'h27010005;
        rContents[20] = 32'h64700000;
        rContents[21] = 32'h04000000;
        rContents[22] = 32'h04000000;
        rContents[23] = 32'h04000000;
        rContents[24] = 32'h04000000;
        rContents[25] = 32'h800FFFED; */
